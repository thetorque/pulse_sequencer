��/  �IUDZ[�d�ޔ���r��,�:vt��S��lo�?	\���j�Y�B��bF�Ơ�K���X<K�X����J���lEu���a��	�=��ϋ���[o�o\;B�p}���˹���	�ҳ�s|r�14:=� ��d�K�A�	ˬB��6W�#�0(�`��o��J����ǡ��H��!��D��e��� l�/���[��	k]=�v���|&]��ё�.��m^;q/��w���x"��D]���^�����UR(5���.D4�X_��{צ�Ϡ�����)Tz���5�lL�$'.E0R�WFi�����H�Y��F����%2d����Y~��ח�4T��'%�Tp�f�Q�an&�eHw/����q�jz]�2��p��hHv��ә��������?9�3���\Q0Tt��hl�F�{x��\7�_x�_=J!�[>�:�+ҩ����J����)��4G�N�|�rg"���Yu�[J�Y�E¿��%�2��Lp��Ο�r0��������Δ>S}?��'roA��}��6��^�y��^H.ˋ�|��HU6�T�]�����>Z��U*f�z�+��eB��i��T(8,�4��(�wM�fJ��Yaib��%OF��N%�^W�Id�A�U�	��x��ݯ�:���v�L>{�2��8��2٧,�s[���m_�{�s��g�ОjR��g��V�=/�>tB��t�R�$Q!Vwc���,b�yj����OPh����==�����?zσV�U/��w�g���E�hM=P�m�סW��k�cԘ�E��wη�L�X(��N�����Ͱ�#�Ìo	�>�YڠR���aJ�ȩ�D�����B�A
׽�`5o��+Ć�`wl��&�(��L��+�済'ޡ)	V�m��8o�����
x�7]�"8�(^_��Pڈ��D����|�V���w!
^��|�
_�����un:�k��T#�s��O՛���J�s>�H�����^�0�^⭧���i�޲0��x�cb:Uc>u�-�W�fj��R�R9�c�vyhH	��AJ��ڶ����3��v��G��}�JO!:�1�B�i(�z�ߏ3}�rJ��ed���?O� @�Bl��Z��D�[n�]_i����ҁ�ͷ���4�a^`��!pO�$�����p�M!�>Fsk�{��Q��vN���
r�fqX��B�q-ŷ�v�٣�'hCGSxW�ky��W�Y�F�e�V93�>��v���h�9$�� ��4��?��E�W��	�Z��y�Q�Қў�Q9ew��������e� /	_��$B��*�IMP}r2|"��b?��{ļ����ꞿ�]�Z�,��%���M�9כ������o�7�o�RW�Lv+�S)Z�ti]�78��@*ݮ+}��{���(h��2��ks�^����(��"P�u�n_�Ӹ ����"$�W����r�O���_�ZTh�>�Xc�=��J�\'�;9+H�A��}�K�4<m����g#�4�a�M�7��B[^f�[��|�Jm飰�4�x�Y�R
M{ ����j��}��F��)���9V\����r��
e\?_�s1�a��>uwGv9g%��$j��)��K�p���<�:����[FM-&����5Q���-����6�1o'WwC��<��àe����xi�؂�I"L(�O$�]8�:5W��]lȖơ�EBG�4�:�t�`Q��!�Sm����
��}��#��;��{|/z�g����>;�0��=X�.�E[d-o��D8l��{�^qm6Qw="/5��q��=���m)ֈ�W���<�HE�!c��i�� �.�"+�lk}� ��뱉��/mVN5nᚭ�����'�m!G~�A�����+A�t�S��ꑟeY��̛�0M�A�ͨ\��5�i3�k"����s�#G ��M'�Ԧ�KO7�$��u���F�����־P�Cp�9�f��\M<�^⑸T��g�qo\w�h�$�I���0FI���e��?'T/x�ȥ*:��l5I�ǝ4;:�.�}�arq
�3�`�����"q��NMLi G�98�Е��������m@�?�����E%e�0��Y1V��:�fU�9ژ�'=A����w
��uB�@�ä�����l�7�哔�5@k���x�q�r�_3�)��Mӱ���v��R��2o�.�ڷA��&ò�$k��b��M�9K�6$��qp���-�5�O`{]k���
#"V�hc��u� �r�|gYω��q�*O(4�]�~����۫�}�[Kng|d��"�M�?��e7{M��:@�	�M������Ov�c�tޥ���$�AԐ��z�@��X��d*ͼ���#�j�k�9�r�m
��S�͑U,���}@����C��p��N%~��b�y����ſ�NI��SA�}��*1�Ne��u�x��$�B����L�
_"T�j�� ũP~�[g�S��t�s[
#,`s�<����T���&� R �����kJ�^��TN A��EPS)�k�IbR�&E�Mc�+�I�c��Ⱦ��܂1[AZ�~��pY��
4��ƹ$��&+Nt,�aSe�8J�襾�
ރ��Vy��x���}���P^��.�Gh�� �@K�}�e�[Aߗ�
���HR.�-�>xwC�<�lmsK�!��/�����&$�_ȔdT�?
]�J�昝wҢԬ�n�!�/�~��C����]����B�� !�s���4�a�V� ���(��c�o��c<Rؒd	����LeڒO��us8�9v}뽏�"�W�;/�	����ǟk�M3Č�x|��	9�Z���4��yZ�+��{�V;��_h��=�IV�RU2�w���ɵȷάl���<_�D�����4�1�@��LVbLHe�m?�?d�24�` �~G�ӷ�S��$��hN��Q8_�
u�4��"8���ݜ>�@����P�̟I@�� �dE�J]^�ؼீ���"2j#�J�7��Fyƽ|7v��i��?����V��`���j)&�a�t�e6���	��j�m�%���j����p�(,H����Wfה䢩C��u�j�rG2��l����; �x���?��'8z5�ט��Ќ�C���S����4�
����P&�2]��4y�`�����#x�#}\�J.�gf�����̵���e�x��Ѣ$�8öw/[/���E�k�"̈�K�$D�vŜk�yJ�+CN[���������TC��O�	̷����WmCU�C�&˲R���]��p8]�{H4>���~Py��S��aA ��Ԝ�jL'u:-���R�+"�D��3�Bs���Y�]$Sd��"�]����1A��	<�6��wfA&#�x���cM���pOr'�@З܊�d�H#+lk��xfH'����G�Zd12�u��D�k��|o�I�;�9'u�vr=?���i� �=�?$7��K<1ا�&�f*A�8������#;.~�f�,���e><YJG��k�[��|QxИ�'��I�����Q!���s�	�7~f��h�A�_ Ń4��ϩZE����j���2����������H��U4ZZ���:b�'�_��垇"?k��܏Lg��z�4`�ަ��W��E�e�`e��G��\\A��H���K����pe	�����9Z�	��!�FGt��a=�m�=�{��+j<���K�4�4�tR&p�C�y
ǥ���<삩'�|���7�)5Ũ`P�����i�~�f�Ńc0.�/���eYh�D*�� ν������+E�"��K�(1��jΨ-�6a	�c�Bm�=nC����>�;�A�bU�7��u��n?5��l��_����u)��1����b:�\�y2:��m���6a��&B�X�VX�h���׮6����w�I62��&�e1}ʑ�3���p*���jnz3��~�ε6[S�쎬i�zx��ڮו��@}��TtZvg�-���dS~<Sb�i�4l˚u]�G��O�S7D�,-���Ǽ��)�_E����"��Mz3�C��!��;?d�Y��ٸ��	l*����AqØ\��3ޙ�g%zz�͖�`�h�g�Yme���)��4L��������
��EԐ�aܬ,�d�,�䅣
&(,�X[;��Zfi�z=�.�}�c|P��(�Z2�R��g���I�Fe�|�:@�]g&���t՝���Ǘ��+���ߵq�&6"�P��P���L�	k꿞��ot��$�5�ɧ,}�+�
��겣S8]��#7Y���\Ε�� ka@e�-�	-r�͑��T�FHڔuQ�
�m�T���L��n2�ز�*8Z�U�^}��+jTR�aX��:d��|_6^��EX����9Py K�!C��*�i;��NHn�ƔV�'H�h p�;�{t�8U�5d�T�	���$3n�*+�wR�l�r��U�?\"�����*k�J����b��,�]"�U����hCX�Ģ�*�xJ�~Hq���A�ojXڍZ�婈\���c�丕����"�ڜzN��
̹e&�5ϻ�]KkH?�V���V 8$4�(�����3�2``��W��䵋��5myB
2bo�����׻�w��5���Q�w�,�3�d�枽 ��*Y��/����9}��Z��n$�㗾]ո�\���뻾ީ�O����	���]EY����3� �����L
���w6��Kǿ�yZ�5@� ��G��s��"�T�p�:6�]o�Fj=�oL�Kt.�p��[�Xu,~$:̾��jU�3[J�i��B��*����Éʔ�E֋cׅ��uOz�V$���o�s^���}�>��aO��s���0J���n��p82�@H��5�It�Z39�~-�LwoM���v�? �,��#�m4���q�	3���kyt��-��B����k��wZ����w��#m�Oj8��{����澀�8��V)c�)y�!����3�b��~r��@��׵W�ko��)���#D}��ɟ}QK��B���:�AN'��%�����ɿ�,^�T����NT��Un�T�Λ��R�Ю��@�O.���?�
�fZ���5U��G�)x!� ��ﰝ1���/��?X\tM�ɿ��`>Wj{�����!g=?�n���ٝ�g�0g#�BIlI�	�^�������7����A��(��x���F͉�9u��Y�Z���tH�>@�ө�lP��f���R�(6Fz.ߊ���V�r;9����A��(��A�h� ֯C<�f��$��������� ���T�3 �+Y!n�7^�]@^���՝��Ecӂ�%*��ޟX����~u���>�rt�4����2��V�ʳ��ո����^1���=.� �7��L$���7H ]�q_��7u�o6xR9d�Q+����S`B$�>ҧ�̐"�l�����j
�	�g�$�$��{Ω���{��r�$}5B�����|[�m�%喿ɦ}�����.��Zlz�~��Sz���%�(G~$�Y^��F��SR�|օ����+Z��c5��}TX��P\�F�~zC���{�i#�,3���M���s�i{�}!�q��C�(/W/G�W2��� bt�|r =�u���.����:!���5�=�א&nA���2*��[(X3B���)�@N�&�J�m�њ\ㆫ��j�׳
F�8.����.�pC;�)����[,�0�Z��B#�b�&�8�*���r�T���&�h��f^w��ǥ�;�ߡ$&R���ºR!�#&�;J���龥t���2���-�l��B�ܧ�E FhN�O��x����t�t��3D$�Ǽ	���������W�!�I��F��M]��W�5��r֭7�\k�Dmڍ�Jb�ߍ���M%dN�?!��_C��i�5d�-7�İ��Z�>U9�y�ȫډakf�܅����(zf#�!CdN���%�6����ޔ8�x#�"��+��!c��@7�����s(P����x�������������\���������_�{%*����~t{���P�L�����&�	�nEq�ӭ�[����ށQ t��' ,w!�"zH�f8/��f�_�~J0D�Q��cOAf%�%�:k�G8��nR�1�q&�����]��S���4J��d��+�h���tKtCp����� H�zI�6$P`�hd.�3�2�救�[�^,C��4��j�1��w��W��<1�.%8ˆ�Ob&�9
�����q�-d�y gcw��иM�+�KT���b������r�ѭj�a�b��fp_ׅ�J0|*����`#���NV!Pl�����0������_�6���r�%G&������hbU(B:#$U��҂T��cy��Q�m�+����tX��(�0Aמ}�S���Y��Jl��P��L+����W3��|\���=��
�1ޭ��GC����p�̆���*�h���Ta�w�d$�,��4�!N�a�n��2�zM��Qe����ߵ匁�EK� UX���i��� ��c�e���%Tq�; X<25봰r�Xت��w��N�f�Frz͚S��7�>ߟ�)N�2���Zq=P��y�8�0�/�n�%��i.�;hkd[{#;�Md�� GְX���^�R�9DZK�%�Bf�H��ua�c��̕��Β�B͚�������y��t�I��'�d�� r�Ăf|+d���BB�'*���*�*��5���o�T�� Pe5a�7�*�mҷ�����<
�� ����R/�y!{\�i��AK�h����̫w��qc(� �V;T�*�XTN�_�{/��|�}�Vg���+�EӔƭO��+�D[���ƪp���y��%Q�c:1�>��,�LZ��I$_Q���'�7�|�8��P�֍�4�U�RP��vO�
�Ԣ��@-����
��B]���WGE���~"��ȽL����դ����\\�m��U�� jF=�>0�i��2ڋ����x5 �˷�bv��1v��'�-�+u���PZ��p�W���U�>ەE���Ug���t2�ʚ��/;������ve�6t�7Ws�\iaNFz���sȑ�+# �Yђ4���ϟE�o�n˓���󇢕y�:�"����Ģ�2B�w�|��c1C����q�PýD�b�c]��F����x��7�1�m ��(R�;Ғ��5�7���<0m�U�-�����C�M5@9������m3�x�t�������R��N�����R�{����bL�=w�?.��l&����ճ�B���?`�￐ ,�m[�H�lA)���m�40̠�<`B9��7� 
�יmK�ݵ�d�l	�7n���B�@QY����;��*��*�Yt@]���A�B����٠���0X�U�*����;b�/z$:���
�(�k���bE�0p�u�m`mV��a���5;�rдDT�z1~���@�ԣ�}���0����qf;��|�V���uR�*�^��V�T�����F�jO��/LÑ��t>Ԙ�����(��p>|h���'s�E��S�4+�Z�)�?�"iNK��
� Vl�&���XA+a���dvr�Ko�Y�6���KSq�;X  ����^z{֯w��]8&V:�����jC=kv�ĉ���6��㐦�u#�`�N���*eN�K�:���+xΌ�x<B5�S�H�W%����EO�x�mr�SJ�I�Rz"�����'�7b��f�{e��'��)d����VT�r�� ��
zz��/c&��,yi��}u�^����_��׃�m����4�xe�4\-��,�Q�eAr��L�a��:@����#�1�����E�@�ߟz�3m���׍߄���<���A-|�6��4u����U6�3x[&�5��*�kL�4w&D~ ��O��Ȱa*MOv��4�x��8e|yx>��!nz�K��2�|��7U����#HBG���n�{��s�a����ry}�"�t���ϊn�)�u��!J6ٱ^T �W�V(Uv|���?5��Q3Mu���Q$�WA����БRv�kRbW�+��C�.�jHH���ս�w(�Zkz�����&&!��"�д_e89��?M��6�5���-!��݁Q��T�M{2�5�[��l_�ɫ�0�"���RFG�����L5�����Y�r�g��=jl������qby�d
,����R��φ5�p��w?��PNQ]yY�p���by��ic���?Uq΀����!c�{����/�-���b����{o�x3���5t�ǔ"^�(~��V���W/���c�൬A��n�8�Zg��X)��F�8��rPmk����QQjR�{�6
�9���zs!�)�0�uK��avW��耕�J=��Τ%���i��F��8p1����m�.u(�X�A��.�:�h�L,�$��]��D��fl�(��rfo��u�t���&�!��|�>��ذ��d� P;I���ځ�)�y���lh����6D��n#�|�Y��Yfn<N}����ÂD¶�7Y��I۶v��H����P�� B�yx�����^���ً��Է)w�͞w��A��҅L�9�/���@H����h�^���V�o��( �c��f_$�_����r��8��������)�9��)'S��O1�,vX�눿w(�cKC@���n��	�,�V�ڻ'Z�~��n�Y%T�9�w�پ�Q�L&�(r�@�h�A~S#��Q/7����e�&׿f�¶}E?�.cL���4����/#n��L�_���,���
�ղ�9;A��+`@�� �~߹u�f�i���������P��Y0xz�#���!� �כ!Oe��&}�\]�� �@���\gas��wI�ᯔͪ��������貧�=
���>�QtE��_��Q�G�v�o0�>^���⅖X��KQ8ܵ`���E��s�TU1�?\����"�]�`��w����/-��vy'@ܷ��!ə�-}@��)��$`�S�ڌr����ۤ�\I:��b���"D�DZv��<��d�`Mkd��z"5}i��3�Q��G����4��Krb�Y75O�q\�(�=Хq�;ܤG1�[�,]�^���}�K���T�~Jި���
2��$�}�ZGe+)>v]?�'���|�����[`Bү���Ҳq�b���&�44��% ��x��� q&�bYS��56u�u���ބ.@���dfr��u7�<��i3�)xM���(ta2T�O�(T��C�(�GlYS����5v~-���zX����Jx��뇺�N��?0rS(��!F���P�ᖷ"�:���8����x��K�m��]s�
D��k�3A��Gx_�nt����(��> �WO��Ue����v�e>��u]�o��]_iIR@J�!��o�I��s��gW)���S�0	�#��NW�'Ѐk�����?}���3�C
l�g8��
�d7�����h��f\Vob������*�72A��f�aTl��J��r�jt�����Zw^�Q8�r�����{Cr��ƽ+�|~��R2��6u��p%��]����!�o�Y �9��b���g�㯛{9"Dg�b�S��c�����e'������7f|���Y�&{GIHUt��8�1�=��W�JC�\?8RqH������[j��@���X�R�0�f3�y�Ա�9�W4Gj��h�rU$�{?��FaiG����:ۍA71p�TM;�
M��'���0���_�1���V�կ�/��yUC�iyk}y�*A����6�C�|�,�#�]���F�g��'����4�?-�0d�#�
⑸ r�1U�~K^��Ea2�l�6��wm��G�!N�*T�����&�V���d˹Vڹ��+�3L��ͮPj$���i�.^�_��\�!��ڻ���5��E�WC"e2Qm>o�h{�;���>����@ϯ#�Tb4�6�kA����2�p�Y�W��3rΔ[��h�(=�=u�J��F����%���P!�>�x^M$��h�wռWu3�P2�$���4�s$r�ٔ`$�i˶a��XąM�<9O�*3�-��S�%�l��;��~ʰ��!�Ȃ�Q���|�4���<�|>��*	��S��;C��Ciz+\�Tw�.���Y��E�͊͞�E���_5�2xjp���R:f߱��3����d�C]T�K`#��q�=6�Y�68"�8{^�&@�w�Ph���; ������\9�F��m틗<���]�^޻8r�N-�\�,e�Ԙ�$1��R=�; �oT}g����k�I�&
S3�;�L�_2їW�I$��P`M�����-���-�Ƥ�U�$W���R+y�����C�rf�����D?��8�P�;�<L�PSѳ�����^���o����-�p.������6y��c}�긂6�i߼�%��Q��{Qr�{�K+�Cy'nMّ#Q�_���;ׄ�LAi�>F1߲��8��A>�h��i���g)�'��q�K"�u��
��0P}���.Ɛ7M�gg��i2��{���X~�4e��?�ŗ+4T0��bml)�?Q��Lt���1�qѨ�隸J�J��G��\�粜֛����jC���ħ0ۍ��íl�&� ��-���%�l�zƠ���;�"T��K�J:��(�WŶ�L"H���B�k�|��`�OE��6Ӄ��F�{�|�N YӘ���@���'J\t�GN�/��W�7�>�����|X �-����w~A�E���D��%L�A�3�0�.Y�P�bɇ�[�V��H�ÙV�����%��:��74L�����*M���F7�jH��9T��@�O�E#�0U�]��dB\�Z3s�M�	)QY��m�� �6�)3��7DkOklr4q��ms���466�#L
ZV%��e}�2![/��s݅79����EM�t_.+$=&+�B�k��"�	��9{<���g�;k���ײ�f#���ۑ�!�j2�,]
�E����̂d�G�م���~��gf���PE�$�"7�+����/h�ș�3�n}^�@�G�}��Q`�V�du�*9�ف����S��hGK*�� ﴚ�\88��4��P�E�2�RA��bl�����66<M�w=x���`AopQ.�y9v8�	4&cr&�����a4�R��R˗!�lL0#Cݜ���͟�cCi��=�0���֣��`��[�r;��~��� ��i1Y�ũ�R9痩�H����z_F��\*&B�w[�4@��F62:Ћ�����P,�;�!˟r����� ��7Ƒ����=�_?�	"�(���p؝��}��2����
bf��`�#��;T����7�7^ūG�d  L�=�8� W�h�uC��5���k�$��X���TrD�Vq�a�����F�fV�X��~�9Ú?}��-�O9%�ᢼ�7��g��^��i^-�����5�C�ن I�|�z��ы+��\_���H��f��f1��0��&�������-�E��o嚊��5̜:���ߧ.�q����.�`�yk9���S��#Z��Jy�B[q�MKV��˫4�A�'�3�;�R��ۙ/��+S��W!���*r��裾��X��^'�!�����)T4�V��3�뱍A�vJ����S�P����Ύ��mW)h���hE� ��M9�#nL�C�ֿ���4&*�!2�ϜuѠ�X�W�@�p�:���iy�u�a�ps�xs<��+8|Zc��vW��>��՛]w|z4���E�H:!��64�فJ�Ԩ�E	�ozڼ;��j�a��Ua$������G��#Z<����!D�p��7S�p�l9c��H�S������f����7e~&��C�T8�h_]������s�/��J�BQ˽�O*�4�XC�m�q��nc}M�ˬ!!�1�=��"J3�5[�t�'@��\��00�.{pVXm�\2�%����L����~LG���5�u��G��d�o�31���*A�eC����l�(�6�]��`ҹ':y���}w�,ŀ$�L�l"��s�P�-��B�|�	��`O�A�WI^/�z�+��g���5�j�S�����<(l?���$x)o�.�g��o����'�@�e���3|W�  +g�;�����_�6���l1Ϯ�g���IH�ň0:�#^]&�V�x�;t��j��
�g�y�������f���{[�hn�A�Ӯ��X��J�	���$b.�LK�y@C݈�f04�U>!>���?��x�L-KA�"��ɖ�1���4z�-���t?��9��W���8�z�q}�t|hf�[�4�fN���u��q��sr�{�{���o�����ߕ_���!ʣ#������tm���H�(�{�0q�V��{)�ƾ��l��CMB�6Q�Ox��'�����X��(��$}Ԃu�n�I:�ŧ��)ugC��R:m����̟���D	Mk�Xbf�0�P2�s	�%�TwQ�;�wm������f��2�6В����:)�N����"���\y���Z�8+R�53QK,����,����4�8�E���{���]�l�P'|E)�d�C�F?���%񀋜��2�[o���A��c�D,
1k*삗��J�b�O������b��0��E6\�7K+c��l�':��>��(��	m�<����4��}/]`��?=�5�I�:m�4����_�$��� .}�G.K�3+.��+Ҡ.�ʥ^�CN.�#a16�@���U[}��s�V)OQ5
eS����~�Y�S<��;?�#��
������I;���Q���� ��P/0�*Dbř��
O5YGhb��ck_�j9�Sѩ�r�SV���'�8>���Q*�M��+�G䘣(X��Pp�/�p�	�O�d���?��J��sρ���������[^�m�*e9��gK��-�ٮU����j���gz�6E�T���s���/�Oњ�+QXV��Nc���-��i�E$!�Cpq1�Cig۞��^K��6 w���?ǉnB���`��*D��������91�9a�PE��u@�S+�0&���ݛ���4�B%�;[�'t���	�9�S W�n7������/x��{�I��YH�X��&o�K\�.��@�������ʅe>콧=���m��G*.�-2�'���"��J���ܪ��a$1-[y��l�_��B5����]�P���~��ce�f!�Y��� �!��!2�XR51Bg�6V	��P�ڷn�t8o,�j䌖C�*I#\�����q����o�h�E{,�M�ϴ��{�V�����k�/����7R}�EBK���[!�c`��g]ӕz��Į��PPl��-kU�v�`����BK.�~�"{p��d�^ҹ0�i���j�0��SaĶC�K-e�/��!|�8�$�$ٜ3�Mr8��(
G���外,��#�J���a9���7�^����xs�&�pO�\w�p��c�8y��@9r�n�����~7ڵ�YG��:����ʮ	�����#[�gm~�T�W�b�	��O"����|�
d��ta�z�MvPI\F ��udcp��\����h��R���t����>p8��h^�	I�m_T�5vV�I-��h��nK�Ac�=�Y3�n��z��� NI{�t��}��+ Xk�B\%��`���E�6#�1�K�XQ�G�̃O^s�# ωC�{�M�����֫K����
֑���*�yխ��Z�˰öP�R�?IsN(����P��(�^�K�ʹ������-kB��.��=��AI-��"e�:��?���;��4}
Ȉg�u\���#��~�yF�B�G��a�^�L����;�Anư��e�+ϭᦲ�($k�r�k��z�V.b���RQUQ�!���Lz�;�t2I]���U�tS����XZ��÷��F��d�>�c0�}�T�9xv�ꞟRD�ʶ�)�<�#��1!#��x�ʒ�����^��Χ�1 ����%%��/��F�\�y�7����Cb�����������)������8 �|%e6뒘�ԃ�їpi(���z'��CfK@I�.ĥ����!G�m��S{pᗅ��y0���6YD3��H>�XG7	�7]�AW"�!kj��������_wɡ0���*O� s+�$Aij��C�Z��/���M�h`�2A+�'1�Ρ�s��I���V]@��&�����3���X H��r.��EuH��"����˖�2ڗ��+�IKS٫�Ʈ�I�%&"�E��gE�)Yezu����6��*.Z�#x������PA���طu��w?���j�U�Y͙��^�`�L��GU��5�q:��0�>�|ӎFeG��??��T�?ۏW���(4�N�!�"8�ǫ��e�T�/��:���-+�9�2F�T֎1}/4�)\m����g�ݧh(�8k�7�Kq0�.5w�sR�=�cl�����sr �s�\��]��[�!��;��)��ʙ��**�<����<e�Ů�zb�8�!��:��fe������wg�� �����
}ߑ�4Z�7���8)&��Q�!�	:YV�_ML �(:/{�6�?p0�L)D\l|�ϔX\����#HH�=� ��w[V�8�&O�b4�#�|#�lVpz�}}'���V<�����`��n�<]�XD��N
-n.Ŧ�u5S������3xB�� 7���
U��uc�)&W�E���F�«�$Z�'����_{�u�r)�4������&��(&!H�E���Ē����
�k��~��ؔ��1���'8f�OSQ�O�9t�*���T�âXV_$�d�p��ФY���ݗ4���QUjՔP��j�RA�"��=���=�Z�p�n�_��G����i6�z\����,���Q
�a��{㯿�Op%��=���2TgI��=�6J����.h������ɠ���wv���/�7{�IY5��Dc���I��"���,��7��oT�>5d̪g.��1���lf�߁�m44.6�7��ܭ�VzKM6��(�	�	�%GBqw�/��z�a��&E�I��ix�a�Cg�����E�)Yr�qԽM5�7�꾓�שwQ�.� ^=���8�.?B�N@�3�'�c��y���'z��mN�o�]B�����^l��]�a�WU=4o�6Hc���8衉Wk9~{CVr
���[���1��7��Uu����&NT
�#{T��;�������B�@ͦ��"�����_�C�k	��nw�<����e�u�-$�N�.H�x�4��{L��Z�֓��`V�TD(���yN J0T���:܊������a
��t���R�����ҟ���ʌ-�k�?�a|�`�1�w�������)�]�-��ݸ�}�Ƥ�"[���K�3�}�W��c��Ҫ�\�� �΁���p�|�rv0_��pV)�p�c��th"O ��<�sx�V*�ޑ�c�2���ў�i�lٶ�w���K2�⬀�Κc7Y�HA��Pi�ptR����%�t���e�U04=8�/>G�X��'��2pV+H��z�U�7_���ݲ?c(n9V�-B�c�s)u&�V�k�y~p'����44�Z<b=����/2�B*t?���@nM��^_:K���b#�������@����v��s���
���i�p�N��>ܘv[�8�O"��I�+��vȏ�-���G�{ZD��[F��*h�;
"�i8������]�?C�I.��3S{��.��<e�j�-&{Câ������M�M/c�š�tj"���=��R��Ч��;G!Ɨ&F:U�&$U���Mʵ���!$C��T0�
٥��mψ�����5�=U�x���#� 0 ���?�&�G5P��L��s�qg�]��09�T+���@M�d��y=<���=��=u�\��d�0� u�@<��8�mQ��8-���f��@�\1zs��;�,'�?N����ON=oD}^B��5m�x���JD&H��t�S�u�c����;�Z��9a8>��L�nf]]����3��<f��-[�������fDb�����$����ơ��C-���[�Z�.��4
��1�?�[�4�:I^[$R9-x�Ck^�ѨZ��wl���d��Tz����~�5���^M�7��yj�<^s���Ȫ���;VeQ�"�w�	�i�瑖�;��#��I��x�S����CZ��������������:�mծ������	�YCe5��u�ӄs��2��[��Q�N0¤N��]���⢧2ʁ"Z
v��yuWj$>=��+A$&7���� i�0۸��Һ��qv��ŜŰ{��l�OAx��Μ�a���gj����I(��<�6�Ãg�\�Qu���F��[���D�E����9�U8�e6�5��sG�P����a�ɢ�� {}猶��a8q?��hyW����C�X.�mEJ���.��ޯ�;��ug���Jׯ��5$��/��vN]Y��D�{��)t$<b��1��WP<q�����0�]a��ج�Ӿ�A��O�äS]s�{���%}�Y�����ʧ�ל��p�������Vy^g�:���Y���\�o���ҬvG��Y�L�c��@�d����%�l���S���Z>._G)W���1�l{l^p!�Vy���2��Gm�����N�X��,Z-�`�NߒJ�I�SXВ��/�ߩJQW��] ٻ-c�3e��ww�쏚Bm��g���h_ �� ?Y�ߧ�6��PnM��w�HJ��KO?�W�
�4p�(=ԈӰ[@h 
b�u|��C}Z?:r���3��v��E�i��~�Ck�	�罸�n0��|���0t���^�:��7Sx����ܷ��_)�1�R�_�+^SY��R�
����8:Q���}=Qk*ݸhwV����EY�p��m��8��
:�l�]�XXSi��%��;��I����0-t�
Ԍ\��߇Ѭr�o
>���Qm��u�ш�YW) 2J���\w��*{�c2�#5"����^�@*MC��<S����N!p��������m7��4h�f%G�Y'u����k���ٳ˚�G�rL�겆+	�lgL.ؽ�C��|�m����H7�z]>��AoL+�����&WI��|��'�������a
?7B}pϨ�J�MI�h��F$�-�p����PB�ʿ���r��>&o���f�'WlƄD�g�O�*�C����H�x��
�+��zJ�>��>%��pS�喾��]��Xҗ��س��4- Uq���w�H����CG[�����ʖP��+�	�C��d������c_;���dμ��C�-}�QfJ����r�5��7�	�h��p����q�$�`濵��"v��p}/h��f���'ZU�uZ
������q
U�i(L���7"��R0H�_��H8���Q�����w,�LL�&Ľ7Nb(��V���1�*�����"�v��	waJ�	���O0(���Q�9G�A�t�q}p���Q~��4F��sh.v���tc����Tn����f�����os��e��?�H��,���e����[DM.P!�"�#�Y:RD+��'�:#��Io#�QxӐȣR�� ��䲩<���m���/F�ϋ%��[ӾM��=�8ͪИz�{*����=7nU��Ty¹'��5�Dk�Z�g���,��Gm3^�,	�J|�g�Qn�ːܱ���R�4�E�USt7꓾$
�Y�`����~�G�����Bp��^2��c����p�4��-m�o�E� :&t�BrH��A1�u���/c�Ï!G`4]�·�/���a:AgN��f:�p1J���J�v����BZ G'�HM����:�n�����,n0?�!��@�I� _c�5��1��ѿ+���jc��G��-M���p��)���{{x�L�MnJ��Wz��)�+�����g��+c8�M�l���@s���u1T�0�2~E兩�?�]/T���M��Ϝ�;F������F,0�oV��d�N�`�}:0x�5M2�ee;�&(}�n�N�����< 9��-�>_��h��.c�|��A��e,���߀͜�便}��kp���0�
��Uz��e��}S�&�)HMVuKrlc�p��#P������녧��-�#R�s��q����/W$�*��C�2Q��,"R��};)���t,��4�%u����U��RX�Km*�Qi��S66��ڿ���d�R��R��q�>&Խ��6��h�w�x�tyM㧘�x}�4��7�bM��CѨ� Uv	�l�k@Qm��D]��?��@<<����4�^6�"�O�U�K	Ƃ�����1$E�['w�W�{�r9H��&^M1�M̈�'J��~���� Κ#��/��F ��P!C�)�t(��:����X���y�g��,�ǩ��˴"uc����dxL�%�2�@!�<@z;s��s�o�.�؏P߇&װiybdV����P� �>yx^�4��yØ聦���(M��=p�����G� /hq͇`��e��s ߴ�wJ� ��N��}�g���	�o i3�������W� #�t>ϔȝؖ�L�z�	�N�����#0������8z�B���号�l'�K�U�'��|�@N��:F�_�0C�(.6�뇽�*��MסP}�1��n�d�1Ӂ;%�cЏ�餀`k$3���+/\	*�����AP!�E��=�-�#u#�a�	2���Vh6�`䌸Zª�֩��wBP4�;?��+�P�weG��
�K�����π�[q�~�@�k%��1�>�S�F8�%Y��3<�W�7��Γo���@�貖9��F�˞m���Z�h1/
;�r�9bY-�9q�zW�D@�����Y>��Q�C5�����MW��K�s.ou˼Cw�ܹ�vŠ��8)&0���dM?��l�-]�6D����H<(�Ө��.$�5��9���S�3�D�GS����j� ��5�,
��UGiK<��"�gɧ���sc�@i2�1̓�J8���i	nZ0���=#�{���je�v<��1�2��s�lh�U�k��'W�M�R
�_Ð�6KMw�C�{%K�WSR�Qv\��Mn�"~2�U��K�y'�@�Җ�z�/ѹ��J�Ɍ)�b%fl�wT-�/�.�(4�x���Xt�C�N0�|r���0��!�E�oY��O�@�'<Z��:���P�X��$Z|Cۛ	>
P�b���Rr� Zs��@��ƛH'x0C!��v�����w��#�[�X"�f��?����o(ڛ�M�X1ʞT\�2�C��S9�
�U��N���N�HRQ�;nI���2�zTi]A�V�c�Ǉ��?�<的J�h�t�Ȼ:��J�fe;K�N��\#��6�g(,�!RuØ��0�����Au�/�m7���o��Y��g�:)+$lԑO|;  $�;�.
��ٌ�^X{UWP0����Y�p`濳����Cd��\i��+T)��?/DO�%��fPqA+ ۣ����ʴN�S�+[Q�{�T��#I(�H�����Ș�^t$-Io�m�'��z��I�mRY�T&:�~�l����V*�f�M~��G_.ʳN�b��G/�T�_�kF}*6\�d:�����u�bz3�݅tҖ"��@\ɿ�-l�
�P᰷�+�v�7��o����fC��y�hz��zr$Y�ْ�k�6��Q1��"����h,ZZ}4mùC��|R����5RDOLK6?���N�{�p~���`��}�=��V6}�g��#�<E����э=�#Wlܡ��C���LL�J��Ζ p�xɘ�3��
�v\�x̀�w��"�Qf��78Z  ���UN�8�$]���@�*��>$��R�K7ܠ=�[@��U�M�s�.�l��4���I��/[���)|A�K�l�h�=�H� �\�g�Ņ>�/��b�7�6��h�q�&���]�Kv�_n�?p����.Q�$����b5��Wa�p���\�1T�ƀu0����� ��H���.E!��\��+��_>(
%�ե�xNf��ouFϴ[�|�<�
�4<��y�|	L�'QO�揲�Pk��S�~}�������"/	Aq.NQ�e�x2�sq�����V1��2���~;G��_0鮂�p�K_ȝxz�S�,{�S�`E��6�+W��0f��k9�i����B}C��r�]69�(>�ɮ��v�ѭ;�*�"��6��Y��� -��޷��5>��Iȁځ	l�S�ZNƉ��O�R���:71�R�_VK/QP�{�2�q�F01�I���iї*#�K�Jp�.l볦i�˧r���_���Q�l'�ص�d�" M-#W lR�����z���HCP���)C�gqr�ꓖ a%�Ƌ������$&�K3~56	��2��z� ��\f_$��C|��)�C�;>!���.�^e�D`��1#}�5nѶ��R�m2�G;O��/��:|�A�92>�L�9�A��#��=�ɓ{�m����ur;�E�ճ���.�a F>z�Ő$�o���Fߙ��g:�r���Л�e��88������n��Pn��^�Y?8��B.T9����;��c�t��lW8����3����M�z��B���,0(�-î���`<,d�6i��B%*}���M��u����h3�&P�ޯ��j�A���&�ƻ�T��!�s�~S	K���WC�k�v�5�q�pa�&:%Ju��C@�q+�t���j��w���Z9+;��SR6�<N�$>��u��k��2�8�=�{m��ؕ��o�b�<�"#N(��8��s'RGg�K����hZ�����?�����߮�MA2{��^������� "�"F����X�}v�y?�>��2#�3L�B����߈��eIh��N"u�<���N�U_�-�nq̒1�"�]Z�����X��7����}��,M����˿�ڥ�t���w!���b'EacW�b�Yy�"X,�t�x� �q�^W�Z���"sX����/�L�=������\��xR��X^��[�Z\~*9 �W�)�sf�7{d��q�d"6���r�Nx�!?���ָB��xi��>%��C��S"玐B�ʏR���9K��Z9\ �P6����7|1���݉^����ڠ��^_i)�،��H�c�i���?y�p1F��� �����P��;V��:��o�!\R!a��M gך:����fM�Y��ך�}�+޺��0�n�s<ek8V�`���8*ǲ��Lp�u���8�as#J_��G�3�<U]�.'�ކ�����fCP�J�Ėi7���l.�r<2.Pw���FT�&ȏ��j?�E/�	<Fڃ�	�x����*i��7�����2<h�/�GʝB��-�#;����4s�:� �b*��I���.r�&�b��R��Z��p�>և�Ϋ����t�nUoNQ��b��4���f�+�q����9���֭	j5�-��#3�.B�f�v*�q��XN&��k��/���i�
��)�$�"��Ac��_�ږA��3覛�+�`	�>���>�X���/��|p�ˣ���9�ƘJ��^oM��ʋ�оV3�2�a������ݨ��}1�O$oR+@x��^掮�n�~�kT�_�s�R�˹jSNk������s*��L�(^Ȩ03��W�_����!��&?q��1$������JCK?�2ʍ�Mabg&M%���\������MI�R��Rj�' ���[lҿ��n��.F�.�A��ۜ;��͸Œ�c�#�S��۹���-ty<3��H5�C}�Z�DH#ce���@?���og�>��M8ji�x{w	;d8d��}`Ay`:��{��0��������V�֊8����z�DKON(.%c��첕���L��똑��	� �����J���v0N��ApU	������A�@Ü� Mpix4~ޜ>e�b��rL!g<G<
��������$��UW% ���g�Δ��T"DR���B����)7J�V	���j,�P�c[�K$-_��P��N�za3J'0�<�\o3	(����$=����֟���C��y����R}�N����/=�q��WHx-�^��(��ω�l�� e�(���m,8�����đ�&���C�4]��W, ��]����|M�@�UUY/,������j���JT�c�4l{¹#�Ӽm�<�}���h�_��&�1;���ܰ'��*c6���n�G'(����!���c����TzR��j��y�'��\'.`@�G库��q�^�^<wY�(��I;Be�|�6a�gL��Y6�yW�-D��9�"�8"7M/ė4cNW�+�ivӸ��6ysO����4�z�m��tl��H��.�̚��k�����g��5BG��$*V�@]y�`�̊+ɩ����=\�|A�V\07�B4;�i�^�=YpqS�o�H�Z{��r��v���'��iɂ3d/�i08�]���S��V��4�?Ev���,o�jX�w�t��i�#�#�<�p�4v�����[���i�3Ne�����p��j��Gb@h�����U�QL&��W�j�ԗh�ec.�%�D(*Rq�o?�AY�a�n���S!�7gn3���XG9r�W���Q�(�nD&\~�7ړ룭���\5��#)`{��_/]�"����'<��FULb<9٥�?����&RD?W��TBt��.������"��3A��r���j>e2�f��y��hV�U}�湋� ��$���x1����
J�".�y���3prO�YQ���i�ܣ^:Nv\y<
G�"I��&� �Uy�pV{�&-w���cL@�������Ȣ���(3����O/g�WoL�al1�۽����2l�A՞^�1%j�(�Þ�/�8���h!��G�|V�}�^��KO���+{�H#���PN�|��\:u6��B�)Υ���s��%h͸��E~�^��"dR�|u9	gZ�m6�-�pcV5���5���dR8�������)���\�2��ob���{���l4���`u�LSR��us�����Hi�֌h;Ԫ�ЀR��p�'v�-�Q������oV�N"-�[9�@��N���_�%𮭝Aqe��
Σ� �i��� �e/��MNdBovQn���4��>bq~�mh�n�;m�Ѐz8��q>�������w��A��)��A�T�ၬASyi���jk�pmH��?�J�"��T���a���X ����HИ��qB㫜����X�}S1պK�%}�Ʉ�4ߓ�%J�hb9簪�kT�:�и�ؚ��yWK-ē*�-�u�h�vNo�E�_�R��7� �Cu%�W�,M!��6�m�/��o�87O�C0��j�g�!���z�h�ִ���{������G�hU���9�7i?�aP��\]|f������&!���#���wD�B=���������q%�oV��
/�b$��؀�ZBb~�}�Hi��@K���Z�je�G�����F���%��%;AhP#F��cR��L%	;dz'��� z��hj#ȴ�Bp6�2T�������U�p��k�,r�lW>Mٵ4�W�`hO�W�/܂����H����>�� AW�E�|��8�>�	���zF��ll�C�<8m���\	yq�,Yq��5B�;�@�9��١b�Z��L4^��8Lp}y9 ��ʨs���鿗�����t�@#c{{��B�-����$aF@��~�[,겐��O�"�����")��J͏���8(*��W�v�>/K�F��u�R�[�#TS��+���kE�0��x��<n-뚻��s~�@�Zb��IY(k�R���^[2����$��D^e���N����g:��̐��ŋ��:4-{	0q��kl
#j6����r ��Kae��ޭ ���I#��?p���,�Vg����3��OvuҤ�?TT| �v�
?���N���f:Y��z�ƃ�"0�^����<�lV&�P�ԘAo�q B� *'Y��s��d���$q���S�w��/�bJ;+�J%�do)����>��U,��V�ü��!�
|�[�گ�=�mle2�/N6_�мxЖ�����V���+�.�#�1ay��Y*#s#��B�S�`��M}�w��thk)���|+�ʿ���7��8!Y�(3~#��	���xW�F;��Ka�sg��Q�v[�=��W�"ǆO\�:�r
��0	��ɳ<��X���`��?�De�E]z����[u�l���<{�9�sw���bf=�|�
�jI�T����6\�;����e��&���{^]p(�v��@D"GƮ:�P� ��h���ʨ�P}�ٚ�� {����7� ��U��	�&�6� 4��J�a;��/T	E$�o 겶Qϻ} �(�6щ�o~��s=w�V��	Q�V���p�N�Xt� �g�rs��{/�p̃��j=���>$��ۃ+����)���@53	�L57������GNݾS��=��+)x73N6->hsp<>���j���?~����6Z8���<��l�	 ����Qdƍ�������K��p��ą�γ��.�A�ESO�b5م%��V��x���r�6;	�H���"��=1N�˿@�"88n\zT�Y����t��=���sU�Ճ��R�X%G,DV��`��~d��"�:��=�ʂ|�p�vݟ��R�ӻw29�|a¹i�щ�g."N�黍��0"�X3ؖ��ClT����\8�EE񘟳��C"=p>Ȣ����BJ�P��2�2�z�s��>Y���M���	[t�zIx/����4p����(�5�G^t>��R�J�~j�*R���w�/_�N�J2�u�����_����/����Y���[��g�SjZ�_��2v�D1R��BV�� _^��3����t*�����Jg��8s2Ԃ	����J&@>��ٞj������4�������^<<|�qk��U�O�"�uىpK73�Uα�Z
^x[]#�|�&<o��|;(�{�f�e|��øa����ڤ�{�t�@S��xƵ_����S(T�h��	�wJ>�"�f�+b~O����%�G��xV�18n1��_���1�(��x�7�kH��f�[C�ҡ�=�}���ed�E�V�+;
���I�Rax� �G�Ш!�̽B�r%��붴/yA8O���E�A�N4M�8]ш~��ِ�@��F<����h�q��=�~џp'�����<�n��v��5�k�-��L��8	v�k�T�(��L�~oy�J3�&kev�"*`T��-:-�/� ˣ�}�eݯ��%̕��@��v��M�6�/�o��-_f�*O3J���;0�g�X1�U��T@múi�Ջ��౅2 �4̽y�f괷j��� ��orNJ�� ��(a�Ł���{�;O�f��]��:�^d�x�:O�`��4�����P���~��%�6o�3Uz~��gH�����(�N�뫌�c�d�[���\��Q|�Pџ����,9���y���:��A�Dy���|s�ܾ�u����~O��5�"k�͉��E!T�n��B�����!�d���_m��"��ڠ]��-j���>��`�O0��E���>��M��Y'TBz��D�*I��?-��Ev���zi�C��<l4���S�'/7��D1pR�> �Qs=�W\�?���2���[�-����<�v"�E 5��nGl� '��+����}훷���� ��ۗE��n��m��L���9MA��j�gR�F���LH�da�x�K~|�3$:�O4s������������(�s&XB��z<i�^d�����V��QK�����Ba�U�t�9k�zj��e�E�'\���+�[���(Q��oU�@�����	�U��O��Vrm#�. p�R4��x�iki����d�sF�)��RD�db���j����p^G�5�Y�s��Q�Y4�-jʘ#�Ѕ=J)��~w�4wݷ�*�D3���f�_\�Sί0��K�;�"ɕ���q̃�wm׃آ���%�\�(��>�n@�=FlY�&��C�㽞�(!�嵓���J��D�/���zW0�U���a��m�S��@�y��sm؝���z���w��N��ڱ\����T�S5�cLDʸց��fQ��Eg����^��ƀ1 ��e��-B~ͬ�*}��.���etK��+ 䰾@!��� rTw��)oLMb~$�a�*��ޖy�2d9U���-
-]>�����v��L˟]�%N0��Ed3e�\�1��Q�}s �bW��������э?��Wu7���̈́����Y��N�G蚤�OJ#�ö�&o��X� q�mޡ5�و�^8��`��9ޑ�iOӌ2�m2,竬#�?����K����bE��Y�_7�>h)��z9�#s��2!f���8Y����Z��p-�ݏ1�M
�o �ҝyɸ~5�8}^��Q�-�;� �k�>u�)4ҕ�wn�~��j�p���E:��c��O���E �i���Q��{� ��Ed��b������a�We�a�e]�=�o��kk��9��4����\���J
���Z�:�Օ3ef^��99�)�R2�S�=!LKa�����Y��3CT�<y���;ľ�L�U��#��HlӋ�@���HH8��I�y������(tW�	�|�M��H������im߹�������>�O��v� �mx��F8�^m�R�2�����S���p���/3VSJ�ϡ�+�R>�o�G��y2T,����4���h��xɖ�b���������.��hs�ZH^-�v[��H\���d� ��|a�7�䶄�24W* ā�vO2���dD�?�}��츔/g�1�6�c	^��Ѐ���{ߪ�_���ϖ�0�3�T{�aXJ���=�	�˩�%���AL;`cT�{	�R*�Y�ن�J'Six�ŏ��E�`���?&��eU���& �Sd�����j�h}H?I2�4s�f�Z�Qܠ�df���]'�l�v��ـz�F1�q�� �Y2qn���˼���~�J�{y[�_�$u`�,Y���義X9�+���kF��gT� ���J}f�����b[�f���9��ps��i�#,`�"��W���@6	��-������rv����M���&��gӏ84P��g�ƪ��R��j�[�x8�)Ӧj{�X����hH���-��U�Sr�B2/1e�y?q:m��x���9e��X�I͏N��cC��dmp6��^�޴R{����{ɖ+[���/�0�Z޳Hӧ��k��ƪ��0�/� ���(-E�hȸ�qb�9�0�,���U_1�e���%;7��Z�{���i�l��������i�����|3�C���7<�K�'X�;�+��O���N��O؟#6�69�&�=9:�J�K�F+�O2�4��Z��3B����TCZ�n��M)������?��I�~�{}Yd�#�%YB�ٶ^����ו�Tj�v�t�Ӿ�7_����_�HYDAi�_�$�������,��H\������K���цb�i�"�=���iM������������Z4����z+ v��2\�Q�x���M��e��L�؈!����LN*r�/�E"�_P�D�m#�v��~�O$#6$S [h�-�+9؄�kz��7w[ �:���;ݔ��E��Űz�J�����YL����� E3� �z=�s	��M��u_T�X*9j�*��4rCAY�G)ҙ8hf�
� ��r犯����B�� f�Ͷ^Ωov2��?�i�]�Jt��
��\�B�������/y٬��}��2��/p/Gv%��N���՝?�ˮp�CG�G� 7*�R�W�<��8䊺���
��g%Ё�o����ֈ�C���^���G��,h?�h�ZX��`/�*�i����婑i�i����3�r^\��y�A���z!n�"b8�*�p��+�7�ϖ4K��2� �u�{�J�A|sAZ�]�|�O��H<J2PZpNhe�S�˷��,�*|�w~�~�І)�_1F���a}�74Y;w��y;��S.��K
��Yc1�)~Q�D��28go���^x���lwqyčY��������Q�XV]y���`����q.����˿�=_�Y��nt}_�_�J�ZJ�y��N�J�]Z� !����U�+"��JJ���߼�	�*i.E��;�m�{H}��]��Gă���� �jq���*I���L$�U�W��v��Q�`:l�����)��vh��n��׊��wO��	�Ok��bh��JH��"������>����f̛�i���}G���|�T[f������R��$��$G��$�G�%��In'wAO<�d�s��<�!qu %�'��~͟ߚrE�]r�.���pk�Z�ڋYƁߤFkӶ�XP���j@0Tb�f��&~��ۗj�t&�AW}g�8�Sg��l�� �l�W��h�萻I��th%a��4�
e_�7�Wo˧���[l5̽ڊ�K �0_�Xp��KY�o��G��pG�.R�7�ʑ�G�h��y���L�1*�GhZDgkޝ+?K����jx��S�M��͟���߅���O� _m����y<�gl���?My�Ѡ ������p�~}YU�vn�T������X�����P�!N���do�I���NZ���U�?G��%?���_��~߉�c+�ro��~-�`�iy�\<ٰ�Y���x03�<�(��`١i����;�>�ez���f��R�Jj�ߧF ?5��Y�0�'�����k�W�U�5UR����ܽ�zx ��Wy��ǡ��$\�������3]�Ց��]��: =q�[7���l1Ķ��17���׃�蠂�=;.�7�jp_6|_j����<�R���
�`{ԋ���C��E�@�a�w�r�g,@�x�K���j���8���;�u�]ҚEq`��;c뒋���=��ْv�sj���bYE$$`����czj5�z��F��u���"�뚐���Z��]�}����A*DN �?�V�bF7�7����M������]e����l�9zD������f�!�~��[����jݲU$0�y�[�����ˊV^���_3G��Бi�[y���T�%���;ݬ�x�
䝩�MGF�m�F5���HB�t&��:C\'���&H9��Bʮ�k9�He�oX�z�W�t���
��h��s���B�D�	(��m��*��e�$����m�1z��%�1�C�N��8�~�Q��K)���kTz�N�s@z �8['��@}��;��	<9pL������|�ʯTK��ѹf`'M#��U�����n��:�J��ڷ�`>QxzSOV�H���5���2������/�ʟ�ȸ�L��!a���^;�LP�0+9Y3�Bfh4�V�{f�1�W�rO��Î����u
��1R�Ñ��4�T�#	����#e�'Z#���r��u�4+�pN�����Zn\���נ���@z��)�6z|'���{.$IJ�0���Z����r'U�h܋�߉TD>���%S��t� ��/7֣ݯ���#��jݥ'�qQע~�����Ω��Y�����f^&�ˣ'2�DW�a�fsց�1��3�I�6��5G}-|H����8�˧¾�$2��N������P
V&:�hV�}v�- �E1.\*+_���\����SuX�Q��8�I�ke�5�\U�f=�����#�q�$����1>~�:;,/2"��cjf/y9=;ŷ��mH�ZP���_w#���9!�9Q���|Qf� �=�~�m!�mD��=��� {ǜ�ｭ�����4�����B,�-J���~��������cM�w�����7�N��m�3�J�c�����F����q�L$��_�@�,�?dh�Z�.�xS�%��v���z� �?g�3ܬǆ����5��f�cIy����1���c�x<r�?۰��$N:v��N���>L�ɵ��fcm	��d��*N��/�+D�we�?�h�>�,��\Eͺ��r���ԃ�&�H�F��}�`��gI�}I�̎zv�g������o!��5���!D�|�(_�G�a܋�9������W̶���� �p�o3#�\	̟_��⌟��j�F����s��j�#��:�b����^�ޫ��|�o�Xo��}�@#�o��-�DR�ټ�O�M��zK3�������j���2:17i���><�T���;�L���&p�]GR�IG� ���b�Xh��f���z_/�S�%B�¦��h�!%2�c�*jo�v����ʰ�:1v�|�r����/�u�͘�R����l�[K$V$�-�EL�s��{ĵ�bt��"M��ĎRE_�n�ji������^!0d�f�P��"��:_���
�Ij���aѓ8aa��D�\o�~{��i\���!O�?U�18G=���� ku��+q��jyX=L��e�"3���J.��(R��^�]���L����DL���=�9��}�1�;��$���KBZ�K��y:rǍ�_A?��\f�R�1�k,�yi:q����6��@09G�dL��4���al�<��#ژIc��xε�$'��&D[�R�F��LԄ��~`R�ǋU���i�/�̃���"i�`�%�[��N]�0��zۋ�g�ݩ�O��;i�Z{i��F6�7��� 5�wC5��y����ah�H��j����AYn���$�a�%A�u.xDY"�������p�y{ 3 ���n<	�\��m�G�D���B<(��*pH�@���k�N.Ю} �ל?�s���/��M&���/'������@:n���ш�p�F��(旇�!bp��9b7�yR,J��<���<��nu@�'��n>����N�R��$��a$�s�Z./�y�t�휭'%u�wR��	9��f?���-1F����)�4Kh�Zu�}����D���1dքF8��e
�%˭x*ܤW1�O��A��R��x��9�u���u��S�q�|��mW �{��Qy~��=�fl��3G��p��f~������*`ч'j������iT���`E]�,-�Z���L��8I^$�x�Il�:t�.{.������L�j��n�&Lk	c|T<@Үp�@pɎ��nvB�b��Jp�����_^��Xkr����2KF,���(��U�:y���h�
V��N�t1Ps�Ķ�����rԺ�"�������Ed�DUj؁!glT~I�r�?�<zDۢ��-�X/�9+�|�p"3���n�S�u�	~h�j��X�Eٝ!c�M">�Wm���x1}$��
nV���D�K����j��/Nh��`8��-�=�j׌�Q�:��J�/xA�8�$�:���ʘ�_�K�h�� u�;��4�^�[��;t�4j��L�-�߬tSٵp�'���?NF����~oU������ԛj4�Bx��ͭ������N|������hIō������0�V����9��S��تݥ��OA5=.����V������xvC�^ϭӈ<FP��i�ʠ�U�W�-��!��9`���[�?�a�8�0q�5�<)7��&�;�����vC��$�"�ˤ"ޞ�&��(91Q�2���e����g녒I-b�=��t6���][�P�x�\�*ݛ���^���J�H���l�qo,F�C$S!-ǘ��h��Y����8�px�T��;q�U��؛&Q_��.M��p�nv��SN���tf�VZ0>��>I��Q�	_8���6��d�����C�QA�l���Ȟl*���!�!��?�98{P���72�o�����#}�D8�L��l63[`�5�ph�a#8�oĊ���:%6Z�0N��7T�~p�����8�b���裧�Ⱦ�1ܧ� �\�'��������,?��1\�dn2*g'i@�e���~��"�\�չM��r�`97Q�z8ʒ�/d��p,�"� >��Bd��嚍{�;Iv�[���)���ٚ���N�z?�S��v��a�˽?:�g��W�oUB-�#�н��/�ܷM�E}���=��8��e �'��>��#Ы$�3������k� �d?��^W��aG!C�3�2H�NMP(�� �?�{t`5eo�G���Pϖ7O�"��Bo�d�I�.@��Wd�b�u�����[Ȁ5���GN���?��Zk����5|��Q?�;Y���j���[C�/�cr5sШ��@S(�Ӵ
{g�QMQy�]V�0~׃�T�G(����pD�� Ѯ���)+�ց9�������
[�zU�0��`��|\J�kR0'�0����m4�jYltƍ��A
�:[�l㏱y�M$�,���� ����yu3p8P�S� �x��U�a �����t�W�$r����g�\+���7���^�z/r����a����li���Ap���(��T�
�S����0�壊��w�_&��;���^rPa�׺����`]ɽ�����M����T�N�Ln	�V8���=r|X7����dX����H�(�f��e�i8���X�^舩�+S�i�--���Có>;<A�=5�I��f�9���e�l�7vֽx>J�����p}l�aʰ���:'���a���I�]9����E[���ݍm։0J���5�"�m�|���ñR/A;dPc�p��zՋ,jT�o�ԓ��U9��Ӏ���S� 6�{��C6`OAx/	�f��)m	w&c��g60�/'����imSy�V�D%%�g{A��1����s��
�U�[���b��p�����B�����^��b�����7�i�E���0*��?~�f��2Qʙ��+�j��x�� �>N�����9���BV�c"���-	�²#����8�/6eo��PK��X�`
t����L{�]/{%y7��~r$fe����*�Rڭx�Y�D���A�_��|���G>��	@�jZ�B�����'�Dz%7�%{NXI�}��a�	8^o�z�B�;�[�3�������䔒��<��]�>�)�Y��v�+K�Pz]B�� 	Srh=�/�,G�EO�Z��0_A��T)2�S�"�kn�WܣN�a�Ԑ�?>�~قz8�?x}�s�7��c;n�y��3p]���wy�`����-�����F��p�@��-[
�4�nq0�u�lV���2�C�W��eFq������&ϚwDk��8���Ve*�����<���!�C�䨋�F�!�y�p���Q��J(O����}T�dHḬ�a�j�x-�}X�9~��m��\��r{j�V�F�;b���2aH���L5��(���p^��̊=��Tv� ͳ,��?�^�t"��䟋���բ�%�vBKu�9`��m�ӆ���?0s,��.Z��5���XA񯄩u+�'�6�Lq����c���Ӡ�I|�]����2v6L���o��a--���E{E���)������a��l��_�B�)�B�X��&~]�PR7�ֱ����zZِ#$1�D`U�������dy�������� K��a�Y�����0�%K{�/�݀�+H;118B>߶'�+��i�����D���h�`qz�vM�3�J5���?� )�!F�W�M8 ͤ��Z(�[G�%$�O�M��H��'�;�_�����n*� ��o�H�9���EL��wFٖ6�������b���:�l=멤�¥+A�ϖ���g�;D���}�7vNQm)�S(NW��l�&o)I5�����&ş��2[��k����g������Z=������Wy�:-�� ��e)]q[�Nž�R:y�t�,����^���8�1�">����f�4�*?[tbm]ur޸�9.O��+�����+���\&2��:-�}dd<����$;�$T��mo^^��T�s�����qL�{�s���{��j����af�e*/�M���z64�oŦ�D�Bj���qf���1ޡ�G�f�]ae�ٛ��Wt{�P���N�ϋ��u�KN����P�w��O2�\�vZ�p����U�y:%'6���J~!/t�_�������i?
�D�#����\�-���M]@�XI�,Tr�۳�=\��RWd��PG�.�e���]+����p��D��Ւ<�#�m�_�oAIR�}�>�%uK�v�.�_\L���T�����	K$S�)��'Y\�&۔Ŷe|J��c�'! �/^\�R����o+�,�bS;664�wҺ7޻~Ċ�v��C��c�>#��swPN�0�I}J�r���P�����w�t0�}��pK��w��Sc��<�ɜ���HLkm�	ތu�@d�2|����/���2��**�u�ܭ��٫�YQ�=��{V���2��(��x妠t�f�s�ڞs�=�Puf��H�K�f�Z	����"tL@��)�Ť1r��ٟ��o�)�k�`%��Ъ㚅rrޣo�x}xP:��XO�2%�?
C�j���a�3���(�Eh���FF��>¤b(~�xE�=���О��7i)h���[��WO�)�� ��┡i����dDf��G��O���ͣ��I�*�����>�h��x�W,���|�/���)Қ��r-�պyk7y�_�o/�H��|�ރ�<�����ī����b�����dւ|�G�s1�M3��G4��ӵ"0n�� (j= ��{�>����S��+�ևԳ��_3>���⭛�*�}O%� �Q�2���OoCF˭�3�n�3e�P޲g�/�Tӑ��~\�$����K�P�X7�v������v<w�w��^��� ��(-��f`S��� �Uq�!o�0��	-9`�?ID�≩M��N��~���9㗮u�)1y�o ����4 ���X��FQw�p���w���� !nmc���biI�%9B]i��bm�g����3�?{(֜���2/wR>���~{���6Y�k�ѫ�;�L�2���]�{��N+1y�?��"	�)�vC�c{����$�,%r�H��u<d�`��Ȥ8��nqه�z��B��(�S}k���r�i��90i��+��UY�s�\ӇCƚW}�[��o�
%��	�!	�Ks�lmg��F���#0D�[]��ZC�8�RW��r�lú���S����3��#-�]�u�5z!ͭ)}x
h��������-�a�N"�����&�	�7Kb>q����l5�bB'��`�C��x���kvc�،���nM�_E&����s=G�����h�� ��\x��H�V�3t��@���Z[pIqoQu��6˯ζ�ΒA9��q��ͼhk�������Fg��ܺ~�<��Cs������V���oaC2AgzK�vkC�_���>���z(o\| (Y�r���T��@��d��f�SJ�	CigT g �UF.��F�k�d��=��T�j`�B���Bh�Do?�a�,�.nѐ����M�\F"�
����@��P'����;��s���:��I>C3fB�Ǟ�;�Kyz��&��Q�3j4�����vS{�1X5�uO�w�Qޮ�<*8��d�o�P�s{&װ��G�	YR����*�k�_�	/��u�����_Q����N��˪l���H�w�ĉ��K��|�wW���a�}q']���� ����G{�w�tB|O��~�����hO�*����Y`��v�w�A?���uv*I�=��~�ojP����-��=`�|��c�ӟH/�����D�&���)7�-Lܪ=�ږ�As�|��L���cb*^�`Jea�	w-Η���j�mT������F��o�S2���ȈX��1�sfyU�5Mq��A��F��ڰş��U��T�#����݃���Ϧ�=�J��]g4�0XO,����<�c1�Ym���ʈ��/c�RT��ܢ�ܑFX�b�@�v�D����k�my��QWny�����s�|��3O��{�%�iS9=�P��0�-��H��}��Hϋ����b�rNS儾�	�Ϡ��<.v~>�5 &,+
*H~8��g�\�ٸ���"x˴n�Hzx��ƭ����jT�z�S
m����ûw<D+˃q>��]��_R�$���!o��;�k�zDa���4�����so��QOG��,ׯ[L�O�sv�NsɅ!��/�y��eg��¼c��8�l �[��l/��K�����N<�	U��4Q����Ьys��3�̨�$�(Ʃ��.j1&��{y��\����l0�j%�v�fC�P��n�ղ|��*���UF��H��G �TI�:���#��	Y�M�{N��hD�0(d�Ĳ��R�l�f�ro}�0��Bg+A�C�L ���?��0�p�F�
�,�Ȃ���+O ��rK�����-ii�Ĩs��҇�?�G��c�g��fdHa����~Y�f�� �xV��BM�l�+q��֎�Gz�(W�:7͏n��w�ɷkT��.�bQ��K|�ʅu6�\��U���2��_�����~��oX7WBK脞�g(<kɭp����1*�[���z�I�{����Ü9�#C�6���֯�@�R!�%O��ʇ�3��`���e�jK��8D���^�0��ϐ��X��f:|o+���; E]�:��EU�zk����ړ2��+��#�vRo
UY?��ay\S��	Ce�#�D�^n�u�$�Q��1 ����]�mi��d�O>�lH\�wj�ه���))�7x�r���G'Ԋ��פ9ä?�au)9q�x�w�E�?�A�sAr:ө�ԟ�9�B9m��}�k�5b���	��)�G�B�/�Q��`�� �-rS��!�# �q���~|�����ĝ��I���<|��-��'�=R�����-�Z�YQ�T�l���u� iTx�A�Y�9�|����CN�ȓ UJ"��lC���U�B�է�!�O(>�}��J�1�(4�����'2��Ѷ�Pݣ��[(�v;�A",K�0��������:e�Q�{�h~��cS������N��lrŖZd}���m:G-q �g�m�y��^W��f�3e�bK�Ђ����E��+l����R(F)/Z��0#�2���ķ�0v�$}-)iD_1<�"J�s���jb�QjyA����	0�P��""]���� �NB��vpOT�2t�� {���$�o�a6w���f��%83Æ����a9�sЫeC���x+��N�
�]���2f
[��M��޺p+�bQ�>}K�n� Xhclr8L6�?��M�\��/�Άs�y�(B'l��lh�}��8%�	���hc���c�L"Q��&�U5��bv�v�r���x&�����%Z9�����-�<|���'��&��Wf�'b�ߍ������n<b�����g��9'�S,��	�?B��-����:��Q���S���0�\��h���ک.sҵ!&�lB�I��[_~�HF%�hIC:y�]���WL5r���E�<��n�l�	�����n�2z��B���B�P�:��o'l�(�	�M<�54��V�lB�uVh����������2��nm���H3�4�@�h��`�HY��^g滼I��"o���f��Qf��s�T���`[���9l�NdH�Ѭ����9� �A{`t�}q�o�U�P�~���z�Ƙ���"f�9J�.��V:�T� ��a��q)b�{h!(�'�����U3�!mC��*�Y�m:+�\�ɛ��ŉ��4�.�\[o��^�b�x��C����&%P@���sb�{f�m��TLa�Qs$�ܝ��BY���T��#������I�'�HT7!X܎�}�ߒ�<�����M��0GB_�4��x���fx�(������lG?����*;���5 S�U�T�m��*6�
�i�zL���Lg��׻�;MA/]R�1���d�h����zr8�����1����;�O~Z��4��A�����n!_��C��m�)n�J2��hC�O��|��E�]yx-�Nf¥�8 k)�c"&jT���w}�?�D�V����*�1mp���i���������M �1��Ǡ�<ҵX��x�x��7�[AV�v{,L�(�7��;����5p)���aC�y
�7�&Yj�0n��e�f���|z�g��L^7l�Pʼ>�\#4U�G	X�L�{IA�{fI�Z�tT\�Y�a-�W��������N�0���Q=!���tʛ+K��nv����H��[p�N�V:�9�GGO[9ć�jG�C��<�"��n�l��n��78�y�w�4�pb0�j�\Rÿ́4�qk�b��#n��?��A �(��F�*fͭ���d�dk�P�f丱���M�[M��w��ˆHoDo�e����N �8�Y�k\d/R���+�<�d���h�E�r�[
��vi���s�M��Zdbl�� @�{,q�`��h�$	dsQB�h�P\��"�^� ��("��X�U�W�gGV�ܶ���G���-�TدI�@�;��D$p� �n���l���M���d5���ύ�OS��X3�ьd%���\�܋ꜟԻ<�Ƙ$�C�f�JP��?�+��f!Ý�hTR�q_t�З�>�]���aN��Ww��+�Y�K����6ekz�	ѹ���s������ݬ0�Ԉ��S���_��IN�c��>����nj�e9���&k��D�ag�5�p�s�F���ג#4]�n�C��\ui����kP�)r��uC]�ՙf�=F�V�X��7�Cvl��|KeC*��	*��(E*���y%8,GP{u)��,_�V^�^��j��Xe���%iw�{��?yC��j���g�V���(���]�إNp5�b)Ze�M�1��d)J�5��d��s~���;ǎG��r=�B�!S�.w=�E�rD!�����܎�x�I&�Cb�X�~�� ��ҝt��\�Q�H0I�����	�`T�r�~��� T�$�.�Ɇ��S��.M�\�OX�u!��P90 ��C�k�6t��nKGV�_��-l�1�	�%G<���ݜt��w'O�6�K�]LՁ0�:���V��*������C��Ǖ�Hy��G���K\_jY%����ڝ�u˩�����q���W-�����ej�5�s�p���h�	���i�R�s���U	Ts�RZu�Y�E+ᵪl\4]��n�f������C���y�q�X����瞒K6͘.]��WU�޷`⢥"�G��+����Lz���1�_nAy���9a �4���OX�,��֖�۾IL����m�Q�x�EGNNyMh=_��P@����
@y��h I�0�v�6��\<���e�����5�#��)[�8�KIv��c-������H�.4���#��$
���Ԣ
���Tw�N}��tR�w��3�	���[�������p����?�dC��}���e�k�������g�2CL!��K��Kǯ�N����x�c*�҄)gK�0Zk������ꨕ��ՆV
[�d�,�WT�H��L'�E��Ͻ���D�[�\\�5o0ܣR=���������!+U�r���T�C^�����\�[��5L�C:l-�
)#�7���+�W9�j[�ͻO�H/-姼���h}*�g��~����t��OE,�}k�C�ƹ�Y99��c$��OE~>�=bE�O�Y���D�{js�`�]���Z ��V%�wChO��t3/����|�=d_:F��·��9�]�2y]������.�_�i�2�:ѐ�(�fvS�����x���*����sO�x�@-�y>�|뇠���y���*�h&��b�7VN�H;z�yl���m�aՆ�l�A�K�ѣ��*o���`�'��s)^-☠��A�����~�6>O�UAW��j��8ԏЃ;J�fr�0W ։2xs���EGI����$a7�:\�83��\}���׆,�:�˕W���F����U�ҿ4Fܠۃ?�RO��6�x>9s���9u��`]�Y�ϭ�wB@���%/�y��ػ$))�|�����>^T�Ωc�[X�)�4\ԓ��������Ƅo�A\�Q�<���-��:u��U�ɶ�Tp]+�f~P�c@�;P��.�~�K���|wޖ�@h�Ӎ(�=�pCYk�hSYV=XA-����.�	��L�q��=ǘ&����ePw��b#���Z�ﯨr�B5eX�܏��J�a l$8�ABy� ��0\U�:l^n\�Md�'��z�Ԃ�<����xg$Vg�!/������B��F���@���`��j)�D�3�TF��-�JRs�.�B��=���N
qDسԄ��Ɨ[�u�8�B <K�(�#�H^��?��S\P��{���o1��m��)�{����V�$�ӮjZ�#Q�����A�{D�.|�@At����9��oZ=3�f �1R��H:K��qBFк�x�z�ML.�-�_�\K�B8wQ��猲�p|��Y,RY�/��vw(Sۛ�l����$�#[Ӝۃt�~��C�^x�3Q�`W�Q���h��-�j��L���&�u~���.&7z����Rl�6�|­?Fd�#��b�c�L��Gb��yɝ�̌m�b��T�
3^%�|(�h>#Awf��ku a�(���d�	5��lnTn��� ؋�H��nC8 O�eCW�Fo��E���`f��I�3�GZ;sA�F1z����Y
�Apq8Nn,�'��x�;�@�Y=T��~�u%p�(�k'%���/	��Z�Mr�p�vr���9E�fq�,I��\R�C��]��m[ɮ[���fg��((��sA�_�ܭ�Ҳ%�VJ @��G�N��=�Z�T#�s�+��%U[�*>���q��حÏ'po=���k�JZ o��f��'�)�f���W��G� ��z������_i��9��&��o&Kye
^�sm�̭��!+b��b�4jn���QeC�.0Ka>�LP�
���t��9��ݝQΦc�Ty3?�����c�'0�?;y�����'>Y�/����j��,�4]�E���2�4��FǶ��!��wx(s��/�C�z&��9�)�����lNU_�c�l���I�h��w �����O�L�i��tr�i�0#vaa�婔��$?���U��k�1�)Z��cs���6j3����iۘ�@��z�E�E��bQ)*]=��6�pxDM��u�I��'�fat �5������z�8��UB�gMJk��r�/SF�p������LM����Z��W䐎�$��eڔ��ɜ�W����5ӱgF~Pl& 9wt�Y�jF��x�=taY�Z�!��3a��g�5�sR�C�rb�&�1����S�uWO�w�T:��?���O.�%�_�[�h�n]�����.�3����֨瞞l��?wn3�I4P�}�䍂��8*s<MY����M"�6yɅޜ6-gt*X
h�o��V6a/kx�9��c[�[��ɤ������bi�.�����;�4������	w���zԕ��N�eH�H䉳Q\Lm���';K�
b�t���������"���-�d:E�8qB�S��/W�dH��5��?����P�� �1v�.v��ߦ��C�B���7 @��#xڍ��3�sp�7#�#�<܈��-8��q�t␄:�J�0i}�	|Z�-N��d�����F?�-i�����z�Xޯ��<��y��A��Kǡ\mY��qŌw�O*],4Kx{B�ݒ��L)�p��ݝ�L����]�$1-��N�eS�xv9x�V&缊�����lY� �3h����H<Xhz�,�n<7K�H���وQ��Z� .�1�Q��q�Te#a+�����VYG��8�o>^�º�YqL�zªAX�
�����O8��]����5λN)qy�u�/�����X�LT�~;��H�"ɳ�m%�Č|i�w0O-����r3�n�}1��%��?*�l�A�0)�n�����r�k�u�q�fpF#���'���KM�kH����%���ؐ��F������g&���8��EM\���pPb�*�)�9*���X%O�-��r<��5S��`��~��+��e5�������c�NEk���vAVW]��X��0��
���V�q���g<r|�m�.1�x^&��<��F�'��0�K���(aeH���(�l^��ȣ����bqh��5;��=8��>�0L��5Q�P����ڶ�V���C8��l�K�����a�N>%�u���SV2%:�(m����V�	4p������m����Zy���Bw������?`.ϐ+��=<?�|Q.�`aҟ�u6�=.T����v|���1��~U�-
��s�¯V �CB@�Z�Ц+�( f\Rؖx[<rD_�7�AS0t��{F]N�ت�p�`Rt+DNr��~�d�ڡ"��dL�G3���f8�t��d��5*lR0M=�x��t_ʹ�5٪�TB;p�U,B��*�5 �ơ
ɫA�L q�X�aҴ��dq]/��������"o%p*v��k��3v��J��_e-b��fK˜�px�#��<�9����%��g�Ҍ(��>������X�чx}/�
���*F4�bo>Au��h��h��2��\9�?�l�.+�O�g^�W�X,����w\S闲"c/xh�\L���lA�+���\u�ӧ����cEk�)G�9�|)"[f��iv�gD6��3�B��ּ{�V��{����7|��T��#�F��V�j�%]K���v̎�\�E�2v4�0�h�����\�&�n�b>@˂OqI�sԑ0 1G��M:�\��\�]�̟�"੽���a�|����C9ɼ�����aב[�+�__��6))>G��m�kqf�bh�������#�#f�n@I?�{Lg��?݉v�q�|h�,9��W�R������D�R|�y��vE� D����O>�1ҽ��ԙOX#�� ���~�P��]譯hJ~��l͡(0Pd&/�0�5kS�=��B�+��Epo>�:Y�w.���nkJ�6P�]@4C�G��eE����)bv@�!�E���+AB�����=��OD�����mfL��5����B<���������ݶ����:����!T+%���%�'�;�J�(��(A��B�06#�bv5��{�TQ�?q��)��ȱo��(�/G�n��j�a�V�$����~F��B��Z2Q���9�a8Λ�|�����2S�	M��t��)_��8�K{�����>B)Ě�^Y)h�
kno#*�}y���`D�
�[瞿��˭n�$h:Cw+�7�]��>�Pu|��_��5�:�V��	���@a�tg6?6�lQ3�:�;�g���V}N�A_{r�B����6m@�%DQ�3WJ˗,�`��2M�|ol�@L9#:a��z&��f=�a�]�t�G(�7 J_�����CK�t�j�2v�+��1�}m��J���Vڣ�P�ÔN�4�PͰ!�"ww�r��[ă�0���r�&
�+mj�~�>� $�˜)le��:�*��%�nJ��̆ԙ�y��=�@�Lt��=nƾ�M�'��,I��?'�Ƞ��B����r�S�!N��n��([�Pd��xp���5�ө<�������kK��%��;d1bRa�W���Rc#,IJJ!��5.! ܯ�1>�F�?��_M4���)�Y�^ ��(a~[\�Wi=���SY�O��G^q!�W_�G�u�����������ڰ�2�'gN��1T9,;�4e��QMk�<�Y�K�5EUTh�z����s��iq�Q���ۍ,M��+k�V���
�=�#_�g�5�1��o�Q���}����<$�͌4�w��>z����S�6�ͷ	,�(g,�O��F�����j�ol���?ʓk6P����8�8q�֔͞PDf]�i?,�Y�[$`(��=�4nk\[����Ȅ�U��I^ph����Eyx�V�Th�<{�9++p���@�1������+�^�2���wL����s����mMv����
~_�lac؆!�_r�C��Y�.��p��@�P/
 v=�(�T� �[���%m�6�u�i��^�)�9��^�T_���Gr��b�Q,*��Ű A�́�~¼Ѷ�#/�y]$}�s�9�����	HԶe+�|��_��'?�#V�҄���͓1`�<ו�Qx"���ש��=�V濫����ZH/FfX~�I�X.�lȦ�HG�0��������v�V�^X@Ru��o�Wⓚ���<��bB�1��vZ��h�, ���[raZ���ߩQp8�$�ڢr������0O]l�C����}Jw1��zzӊ�X�ľf�㻿`� t���*O�xٷ��F�D��#��'����$h���8�Q�/il�+��#����Ք���䛧*��*i��q������F�5��E��N-10�өi��3s�7�Ŏ܂ ��K�˞n�Sļ���|��6�ݳ��H�-��A�1��B+�Ʉ�;��c�/"6�
o�:Y��;��K�x�}�A�;�U�SLyM�QTn�.Rp
��"f�Kl��gk'�8m�8ב� �Z���p����^r�H���`>�2<����T�����,��:|ZR���ڲ�2�]=��H�qX�"5�K���߽}r"����w��J���o��l@����ibt�s��j?�E�י��-J'��('/�@Wj��EO��4�o��I�]�v�%���u��8������{�݀O���Vӟ��Э��=��gyEL�>���K�r�D	uc,�`ɇzk�V-�Y���{��O�ܒKS�c��E8g�;G�ĝ(��GӼi�ə��� �V�%oz��Ϟ�СʍK������=�q�e-mo[z.��?O�N;৛��ۑkJ����e�zCG
�<��e��g���x6 ֙��l,R�[���Ч��х��?V�.��D��sF�?>l_gM��̔�����_��Q�� ��w����P�$��VYa8�x���=����D�}��x�`��N����;NI�����2"]frp|�}r�S.iJ�xNs�S&��v7l�i��v��]��}�:�Z�"�jw�Ͻ3mnw�*j�Vo��%�B�LZ��&�-#�xYj����Vs�U&��'m��bRχ<@g�����	��j=���$ .��IDuE(���?��b�92_� z����w����>�" �O���������8�7	[�����f�����}�7M�Fht��/�� I�(����:^6K����Yt(M%�R/䆽[��0��H���'!]��?4����1��'^�;��M�H�"�]IE�ی>�;�~�1��"���F�k���0��(���1�?f�_3V@�
�������z8ˈ!�&��+����)�7���M`���(�yK2'q�er�Y`n�F��X7;�K��\��'�K�Z�bm�e�x[��M��	�N�=�n�����:�^���|h�:=��nC3��r��U�GX]ql�w�1Q����M2��B��Lh%-���-�R_�e[�>���X��졿P�$���Z�g�#
�?n�79�9�(�+4[�UF)Bm���k5�1ag�cp̪�K��.3��,:��Y�V��� �Dl��A���LE~֖�����[���Վ��u�(cHFi��MK~>�~8����)��Ͱ��+l�"]�$}Wע��5)�n���Ҁ[��=�Qy^؎��h�z���<�R6Z� =����W*B�����%fՈ0<�G�m&�M�0	iF��c��֦	��Xcٗ.&Hhi)[��%�i�[�K��]����B�m6檐�������?�|�M��.�u�`s[P[�zY�_�D��:�S"���q������)�F(��E�`��.Y�#Pn8�JJc|.�ؔg��Zo$\E�Nʘ�!�f�Ao˧R4�������'���6x
tU׏8��V�k����v2�� �m�ȩ��HMS���ԌüZ~����^g�e�+�Z����ɣ�Q�#䚠�7/mܖ�-_���=�av୿��+��V�m}�����'��5YM��jK8�K'��#Mrۼ�~<W��f �lL�mc$ea�y�c�d{�Dڶ��}��~qf)Ȩ��W����&�3F�P<#������=���.?r	4��gh}$��"�7Q>�!z�Ef;X"Ԏ�OH�N߃�f��?#q��&�HԞ�Pն��^�٫O�A���Aj5�pɮ�L�Q*����rz�\jg��v��}�W�c'%cc	������0W��]
5l�W�0,��1ʴ���b	�RZɤVM��>��*���p�9Z	j��(<ʽjm<uV��uAhy�B�<�A�	
��/.2%ɭ_��G�\��Uf �21�v��@�	������)���ق��y�>� '�-�&K�I���I�D��,w�K<��?52 1�{�􅒽z�®)0�S�&U�b�q�H��WZ��ϵ�
�0�˦���3��2rj��Si1l��[x}U�����Ě��d�T�����Nb��Rd���y���07k�5�bb6T���dZM�E�F}��F�vzQ�ہ}�TSw����ys��҅��="�j�*�|��dZ�S	���J;$aX�Vyn(m*x���#�q *�~T��%����Ž�2���>�#�pu})Hl" y�_�/��p�{	��P�ꣻ����$�-��{ږM�Ik��F��]x�E4.[1�H�7��k-��;���j��s�Xŭ�lk�yz&ag�&���v�& XH�>0�6��A���x�k���t63���x�J���A��h7�a�v%JC*σh;��\�ě�կcC���R�ǜ]U"��._��҃�9��P��>��P��R'Kf�#+a����`�ԓ�`�rM؍��������'�Q���m0Y.Rd@5C����Q����g�Cv�{NRcnx��/ã�"6��o?�Y4L⩅bV�s�����hҜ�������?�ణ�0i�!��i�J=�2�gO���zϧ�&��:��C7�U�d-׽��NN��啖*b�;.M�6�?V��TΆ���DV5���T1��N+��Ӣ��@uZ��)�1�16!�n��3���'���	�qx����s���r�~򥟍�.6�j�JY�R�F0��5s�m��%}����y���-sL&n�<?�!%�V�؈̅�F'�4e�����cFU��>L-�_�8u	K����Vh^އxr����̡ߖ�BE��Ԙ�a��+�|��ݪ���`�L��J�<G$�r�6#���ܶ�r�����V��W(ۋ���� �/9@��Yܧ��fD��4M��w.�0\��(��p~�$� V�C4�6�>��VJ��!�O|�ORԓ��B�p�i8��h�Y=
�a�j%�D>�'�oQ��v��N?�V����J(��ٮ�I�Q~���� S�T�Dem)�^��bnV'syE���Y���2)�����؜��S�&�����1Y�Z�>뜕d졌5��!���v	�Lj�II �{�w�-��`SI?�l��(�V:<ʯ���A�-.��ޠ�w�N��Ħ|�}�ԝ֑��a��f�2q�p�~�cGM��9s�ɛʃ+d�N$oMSa��t-�$~��>1�M ��pH"[t���*��F:n��+�f��$'>�>ڼK�P�~o=����0��K���E+�G(��
�!�*���I99��X�K0�Χo%�jG���*d��9u�0�,�W/>u6E�ߝi(�{� `�.)��Y�A�3�qX�*z�DH�Sc�����@`�p��p�i���C�Z
i�X�zrb�L���l�V�!�'���amoa��L�Ļ0IE��i"�^���ۄA��ׁ@W�֎9IAo��L�Y��ye�����x��@��{z��<h��IFW3i��]�/S�/�=ynV�ШƎlPY`�����s�x�����&��z�}Uv�����˷���|�yE�q�����(�T	Ҙ5��;L��� A�� `�=�Z���f�<W1~>x�����1D�w�}�~��vh��wb��c�c�9�y��@š�Ob1H�`�&}��l�{���S���z�����V�i���7mʬЖ���b]�}ݴ��
�{�h	x4�����{$�iy���	�����/�U&Fk���HʇPFN2�/��j���M�9
�֙�,�u���?6�ؒmi�♻U�bv}�K��y0�$g�_�%_�'�*&�������o��I9�O�������<�5�s�z���$�W'0�� �ϠmW��������0��64�z}&փ�_P�Ŵ)u8�'��W6�yŇ��(���\�Zp��>SM��#��	��.�w%�i13�V7��
T=��wB��g�e�!uW֛�����
�lbK�Z�%q���������@�(�J&G���H�O�)(�Lm:�X(�5oBr�%be}�2S��{�m%@�s��12��J{=�)U�BK/�G��{��+2a��� R��W�|�+Dm?'�#�������M��-��`�#u-9���/�K1Lp-K���>4O�q��(�ɸ�����3rOW��Ɖ@�?8�����@�����wKp��u�i.ho�wg�7�������Q7/&K�*t���k�h�]��ş��
`#:T����7��Hw��`�E��u�&
��"�0��^�Bg�lR~,M�l'8C��#+X��Bv����?'�X�C����lt⎶C+�S�֔�N�ȿ�
{K9���}�%��I�,Z	a4��{�n�����k��c�=��˧�8Ot BVE�� �3(��ҁ�i��;5�o��H؆M""���d��Q��-�Æ-�T]-���N6�m��O�VL��XĠwW��[G,Gh2�*��%ўv�/Fs�~�Gc��s_,w~��{�6��3k�t�Kt]�"13�Ʉf������V�yݑP"f�B���^�����\�/$$���t,�"5�I��%/�۠�)H����;}�R��Ǔ����91�ۢ�IU��Z��.��4c��*��*0����0[�I�i8f�O ����S���%�o�y�nT�@�Z�z�& �Z�~c�f�����]�Ly&�w��)�Ö�E;�`mh�u���s0�ƫ�ܝHKcKNw-�� �x!\Z���kk&'���,��/-O�*�0ڪ�K�!��/�%�0��NR�%���i�XC=�ߠ
�uu��,b;�aA�Qܼ�ա�&~�f2�N�ۮ��8��=�R��ޑ|�1���d#%�����Aʹv�ʇ���j`��D�)D
�.�JMF��R��&�$!lwӍ�e�؏��-p��O"2���	�6U��:���hl��L~��*�ӧ�K2���{��yn�r�Uv�R�>��x�^@ka�]�u��xvz�m�_F��SWM2����g��漒�a]ꃔmjs,@�>��"Эcf�wRw���=�TL4zw����~�d:<�K�gUV�٠�����(��|Z��
��Φ��l��Uy���"��Tc�)��uE��r�	�2��J�m^��t��G�����/d*FD�&u^~0-_'K�D�S��r!gS������u�.L��������Kɋ0YǞ��!�K����MD�x��cW�d���fO�r^�la�)]T=��U��?qB�e��*�6���"�y���J�
��E�4��ν�s
��²�������i��"���
�bH��Hd�h����գ���ml>��4�Bl4$���	�6��{jw2�h`��j����~���b_��T���f����n�o!�(c��$����'�S�<��|t��<3��۟��a��X�ԍ���5��z�=��lG`��r8|���2�/@���.g��s�~�,�;R1k1����{�u�8�� 6�(���/r�kɇ..�`p�T�K(���A��;d1Q������=��V4�)��X{5��4Es|��+�ܼ���(D��Ǎ6���E(��a�;�&]���-��Z:ջ��h�[o�^�����$�U��;��G�c�2�%ˆ�X��ŝ�S���e���qv�@�Dgq50�oLw����hpOHE�"��Q��;j`����Pkj]�C����]�"2���sdQ��n����G=k��VR4	���6fb�y˹�}��R=ס"��,\d�J,����6A�,@�ښ"v��ȗ��TiM�=��~FR�'��.���S�!������l�y�_ju>�j�Σ�,K����Y��M�ĭ���a{���m�ϓU�v��.���G�Ұ�Ȳ7����r8�`�0@�wຼ�V�j����_:Ȼ���3�K������U��dJ`�=d�l����{u���ߞ�����~3 h~���J�#ig��i�Y��|��p�ui��`@K@:6��R�V��D���y���ɊM����ț�e �$ovSSޱ>�����s�eć���
�K#����������9m<��וA{�&����L��R��L��鐷o�g�,{�a8����Tc��X�_��A����Gf���9�
�#:��P�����a>8�[ 9�B�l�V��V��-����ÛK���#,���&�~X�J�Y��Kd���@m�݋Ň,�THk�H��`FY_-�XI���,&�L���a�{?i厐���~�n���Kԁ��բ܂�m��(�A5�	�&�,Ȯ�y��Wua�U�@�1e���wė�/;��{0g�]j����jc�_�-��5ɛ�E���ɶ#5�J��h����؎5���l��0���j���ue|*߬�u���a�!#�ȩ��."�[�Lf=q��g����q�Ԯ}�|�K�+�9@W*�,��/J���ڇ�)�V$ e����z�dh�G�W�2�[i���M�A[LCf�Udׄ#u)�C��V^�κo�%�>4Q�x��٩��tJ���$��q9�$��ϕ�T���p�EW-����[����$ep	�7��L���0yJ��
O���j�J,�0�5��|���Ӛ)�ϓ'uF2���r���T
�u�99��3I��x@l2���z%�P$Z�S�b�v�Ȧα۫�eXV���}�՗����5�bj�}I\ҎPw��}&�x͆͆O)�<!��m2I)\�������/
,D��RC��ܪ��-��	��k�\��sN*f�]�Z���I��~�$AW�������g��?������Gk�&�r�u�.p�а.=���ZW�_����s��k�C�.Xwղ�3q���+8a�&�󩞁���z���ǚS���H��>���y��(��`*��G��\
Q}��,�Ϡ��Y���~��(�Z1����`"1]핱ymf+K=�nR�ls1I_���c�� ?ǥ��?��fNZ�i�;�2��"٫�?��(H����SN�*Q5�\?_G��u����L��}��M|�K��o[@��k�5J�h�̺%M��bᬝFE�����R�$��-�����j><�BG:W��w�������׽���=�8m�Z���I��-�V��B:�Ad�t�k�H=H���p��m������K%Nn�e�����EaD����2c����iYs��`D�sEW�����,p
�W����eHz�@��z^s������Qx�����B7�Y�V��2��N�C#m/c��e�F1gj����vɗ~��}�o�O�ũÈߟ�gL2�N6�.o]�eKF�/��mM����(wxć �mT8�+2JW�n^�ݢt��2��:~�Q\�g�(���^cG�����_bPL����K�K� �����D��P�g�\zC5�0��������8� 8h������v�Kc_�_�0ʰt[�A��*�ߍO�k���>[�&�4�F���Z�Xc�%̹��j׀h� h&76{��C>B��q~�T?�&M(s�a���Y�1�F�^�?S��:K:`�4�ő�>�u��i���#����	lL��<(��1�I٤(�t��ۧH�5v��J��Xt=��j$�#CK���y%K�[��M<������42�[|P��W������ӯ aB������}��ߚZ�O�*��0�/�Y�r�. E���m�͛±
���UV��h���xi�gn>ժ8�t\��;�G��gE0�8rn��s�<IK�+��p_�B!��n'R��e��������y�(�g��>+�R���6����$���Ǟi��:ۆ_��&���-��Ot��D_��<h�y��Y�=fr5lI����TX�1���O�:Կ����r�"�V�A%��[b<��*` ��V��mu���
z^��Emۤ��̨ӑ:�%5�G��F��T�9g2����^
��˖2��g�ɫ����r�!��-��1{�-��& �m��ˎ&�/ ���&/�#;�k��j�:�k���ͽ��]�J�g��P�(s��ڀsdn��Z��A�Y���%[�ў0[��]�iEB���Qf�/�,�NXc��1�V��T��[�
z��tgaQ�vi�!����F*S�y��I�_�=�7�����yi�"��
2f`$@|c���A�g��S��W0���,��z�ni�ϭh�W��HBqEiuc�A���0�P\��q���	b�$'�/�� Bl�����}_��t5<����V��J��̷� ���2�*�?�9+QB�zT]�9Re`��)��sV*�ί�k:��L�`
���*D�,��Q�������oThK�����<�YLS�yL�d�A9��f4`�Z�D��d}���A��4�Ю��8���n���*'�{�0
��[i��勛W8���c0���b5�����;��d$���zp<�#�V�$^l�6u�~�8]�B�t��O�^K0#���D��["�����hL�HfZ�ԛ-�:���v E]�(,�j��8Hk�^$d����ƀ*8�q��� ��
���_�-�n�Y���Pr��]�R"�\
6Z}J#��Ʋ&��YG(� )���Q����4���Ic�������J��m�2Æ�񈄶��☌����e��`)-�1��M��;�B��jR�/�/�D��y���ڇM(��w�5�"�+��;-�٫B0���_�W��!�^x����	Qya��|��Ѡ�)]���~��k	gz]�������ݰB��������k��{�y���	ɉ\�`B�H�0��?��-�۽g\�$ԩ�}3�@vx��e��#��R�v�J�Qk9�L�5��)���Ri#��xCU����*����WbN�87x�ˈ���3)_��ώx�9``��Uޞ`�Mi=�s�&�e���;���y�V<�5@?�zV�on�,B8��H���>�$d�/����EB0��}C�����>�C��^�j�_EDN-��BDC� ��]�x˶71�{}��Yc�`z����ǣpd�r��o��H>��!}g��~��L��f����E�;4g��Rݭ,02��!g�:�2��C�s������\�͡�*1���?��VIyC\V�I�2p�])H�i�	�*>gs01s[�}f�A+��3� �0���TS���|	<6cS;��~8��>��Ȉ�	7�|V�e^�x�;ח[��䗩eù���ƚ>z����ŀ��2�i0ΰ�=�C�u�
�6k���49�ax��إd� Ҁ��X���+D@�w��{
݂���|�^�l&�O	^ �U��i���/��q�����@�wU���#+�G�C�f>�l~�(��O�Q��z^p{9J��Ts���]��o�uuy���<Hp4�i���vd��_��G6��7k�M˻[��;�ȵ���G���@����!Y�ӿ��(�  �l-Tڴ�G�i�0����B��_l�"��hV��#5N#��N'��FɵPNN��"�I܄k�D��g%�B����A�Тc8$__�I�p���p�̅,������5>��E����{��ɆR`V�QF7��Z=�W��P�Fj�~vF��)Zn�Oz�0v�Q��W����O���Q~�y���1������(�Դ4�S:�by�j�L�3|}��C�RC����悴�f�s��K[?Y~$��Y�h,��F�i�^��pk��}��8�(��Yj5sMZ� ���htL��`8GT͆�P���m�2��<��8l4���7J�^$\� ]i5�OӍ�(��0}�A��RD�|C)L����K��&f;˗gL
7��֜R�! FM<cـ�2~� n��b�]�_��%�>.����zS/R?r��S�&�~���Ȅ-2�P�Nygk���O'����B�KإuC�#E��ucƤ�m�T�6�'�0���������0G��Y?�[C&_�ߋ5����*i����媧+�~��L����S^[׊��n-����U�"��������)��ӣ_��+��{;�~�E����kb��cu�Ħ.�D�PT#V��
��d.&�]
�E+���>,�J {�v'HX1@qI�����F���C�"i,(��9��a�R�}��=�A�R0�'hH- �
��n�C�0P	o������B�8�d����J^���-UT��o��$�:���Y]����TՃ�0^`�Q=-���<x�1d���w�V-˽�w3#�x�k��E�� <�&�<O�O:\b�x���� �գ�\�d'���u�&�p?�}i�@w�w�uCLB���)��UEXAЪ���g䌙�tj���ļ��Tk|��3�N�<��"�8�9䫺��������d��v��0�1��P��,�*��������C�a�Z{x�Kr����u��X��f�њ�T^�+�
b`ښ�K��y#8k�+��e񆶨�W�������|�(;[o��7dOg-���*d����&�4B�d�~�z
S����W@����`fv�9�b�<kj�����Qײ��hI��45E߯�����w^}@����~�De�4wy�*���֜�)<\/{��.���D�����ġT)N6���HM}x�Y�v��(TĊ�M-c�����)��Y��LwIk����)%k��G�!^����)
�]}��	k=��%,^Q�H��>�"AQ`�p|��7v�qV����vƜ���2&���^I��#?"�4j��bc�=�X[0�ӑ�g�$�*:`Jl^?'
��0�qzZ�C�*"�"��
4T%ٹ�]���P}��P�/��]��ߟU�)>��`9�R�M�=�\�!=W�6��̼�`�9���,HST�QeJ�O2l�G6\���c�?�0��oN�e����T[B��*�jZZ�B@�vp���sμ������U�}�bjl�_�974�5�Ņ��K�79�ʤ�ʴ�߳�PR�����(�թ������A$HM.O${�x����E�5$C��	�`�ИMjIJ��0�8�sy{�%���3"��<����.�h���fM>��<\K�����K/���l
�04����wEf/�Hy5�{ék��2�y3��`|�$�3��m�#�X�3~Ν0z�f�{A�!��+1fVA{6(�>ȥ���`�������=�XI�l;?0i��{��p,�k��R@f��	�+}����X'ϵ��g��q0�C`v�&��[��2�H�9w+��C���d�D1��S����ҍ��������`A�,��[��������>�#w�����o4V�ob�,I�4�GSf�뤂J��Q#��ƹ6e�����K�:K�s�x��J1Y�翄 ��/:Np�1��L���.9e��
�ZEp�fg�)�-jJ;m��I/��̧W!r\�Y�R ��[Y!^����L��$o�k���˱����m"}3?�H�>��Eu�|�Llt��>| ��h��X����5���>n�a�#�,e�ttjO/�Q��,�1k����;�;����w?�m�KO�^uW���we)�����l���� ����V9��,sO�yrĈ��jw���E�Y67~�6�ә6����1"A�%�JAye�^�x�"p�V���L ��S�d�W��)�Ъ�#�m����Jk��&�ћl���Ɯ
��!OF���!�C�SSƄ��0|�_^W?7j���^�)B4*�x'�I/p �GQ�.�"p.%n>Q:�9�w��`��='cu߲"�խ,	 {.��Q��G�7��k��Zx�Y��u�Ɗ�!�G��.ޙ�[[���)��:w&�;5�b@�i �N�߽�q	P/rY���&%���� ���J�\�����"�8��y"�T;4bX
����'�s o��R�,��n��tR�/��`	��o��iK�-�m<�w�)�)��9���N������?�,�<T������D9�B �����db6��_����N�-��
J�A��RJ2¥&���5���I�{��E]f��P�ZE$�L_l�q�J���� I��Ԉ��w6����'!��Hf��>E�����?������g�ϟx�����%P5�J�����*��d����o�MPm�:��CCB��ѝHwa�i��I��5�D/�¾�����#=�g��y�y���[M��2Cz�K̺UgX[0)�I��� ��yy��كt��}�'�~�p�w�y�C-�*-�Co�K�|[a�����n	X$>[��0EA��@��5��EZ�"���np��H/$�k�{+?B0��us2|u�W4v�����u?xE6�!f�xn|��lg��c	+��������5巐4��S�=^M�	5T�k˺�K>q�k�e�5�T����&%5Z�#0Q�5{q`N@������G@d��B��.U.t�2~c�����<\�y�Γb�NBQg�$3f��>aA=_$��V�̷��rsc2�;b5�Ś�����(7Rcf�L��+���Ec���Ƚ{�f�m�j$;:�E���F��Y�pщv����X�}j��P�&Q6�*Wh.���U��@א��)0 �:�؝Т��Z�&>�g�4�w}|	�O�v�.�g�O���CBd�@R��0L�q�ZAq��-BLg��*�b&r�]zm��to�r3����0NQIU�ZMf�c��UnJ�!P���U��9�߰��u- X�,�xB!7���9�Tڬ d�ٖ�lF|[ .�?�&N�$
������%���o�	�a�qG<��;�����&u�+G����G���\�+�3��g��x<o��*��7�!+�>X������K�9*�H?��QG����~�Q7	=�Q��
j����t�3�D`j����������h@����G|`DY�$� �Wd��|��u�x�e�i�Ӈ)�"~�"���;��#��-���0��4j@|�Q�3:�K<��ܔ����N�g^�������<y}���/c�[���Zrz$=9z�j��j�(IC��ۭ������{B�U��Oԑ�_�)�)��}%����陫Ԓ��V����<�j`��s��	0��@��.�Bu�EQ������6+@���7��QLf�g#rܻխi�镅qԤ�xVh���\��K\�AV����E�?G�n-[5�ڟq��u�K�������c�5�p�&_�r�ǫ�v�
�*Ɓ�(��p)��MB���N����}�k=A^�ր)$9)�;�H�>�
x�m"�%��+��%W"����Q���
�U+$b�1+��K`g�m�?�m�m'���5�G��!/���J�q:�G���i�D�h}P��ΉTG�fПr��-laz� �|����44�'>��m�����4�T���H�nNڢ3�B����Q]0z��{_�]������I�G8*a��v�7{�nr�i:�5ŭj���2{���js���[�C���+��}5w����� FaO�W:��n�R7�DOL��|�tЦb���W��8��K%���m����a��vX-��oi�O ���@V�9â��<�Γ�B�D��S�*�S8tƷ��w�҉���ŭ��Ї�貇���<a�����z���{����P!���T��?���W�K��B���B��"����B�Ҍ�g�E �x��5�z��%�a�Xp���p��d^H�g'[�zoawe�#b&�r ����1j�]�,��`l�j{9���b�*�����=J�M`_��L9����h��<U�x'ߜNjbU+?���r	�}N�>�����v�BP3\�M�	9F?◐ �!�#n�U���G�Z���*tgT��\���VӋ��~���^�OН�7�%JN�*���m��5�z���Nb��C80/�k�lݙ#V�2�7��,ժhm,���fil7�o"o3��P�� d6���P+x�:��H�y�}k���:�"`�B�#oT8����b�-&�Gk>���}v�D� ]��XV(����7\T���s�ퟂ�H���]�M��`V&w����b����ڝCLZH�"������-�Z��O�2E���p ��	"<\��PUUt�A�	�q/Iw�~���`��X��Ҩ?�@<Ɍ���uJ�M[��R'��������p����?l����"$"��J�j���*�݁�������<���
��
�Dm��=8m|Un�����UBv��ti6��-]��Lʼ�7��^�9iX��R�0D�9E�z��	��,�S�T���xt�T��WE5|�G
�t`Du�`�����ګ:4���R�J*�����X��G�uf�vGC5�U���r�� q���~aP���O��x`����M�����?��z�����t�xS7C�g��`��
�@}������+,�i�T��b_u����%�2�~�\Ex�[3�E�۴O~=ǐ��I��F'�~�E�R&�)g�L������Ar�1Yr�L6�ݼ�?��#����6g��3O;�2��4�0/@�LJ�<i{���>�h�qA��L��{�{l 0�h������L5ҘD�D!9�YrS~�H9�N�RT7�+RE{@0@�{qw���u8�K~�ڷ��p�����劷w����A�:��\g�*ڡ��NK㚴�t����v���S~TK96J9KA��#��]���^Ư7k�)��A�Z*�E@)�$`>�<��9����9�g[���a�4C��� �{�Wm*�1���<�nT]�Z�����[���M�Ew�m �S��ZU�3��@;�?�C����=Y�-%� ��Tx�]N�'Ԡ�"�v��h�g�q����Gl��t��R��xwB�;:�������y�j҈�C������{JE@�|��ʅFy^�� ��;��0(�Tbk:���_�������G�w����@���"�Q��F�,�r.�k©m�I�jL��P�}]aL����VISs��eL	>�@�K�]���jqk��:� �7���鹊�m���]�S�`)$A[[�D��>Sק��Z�o.+D��9����?e1����<�H$��]AR���J9Bѷ��s�n��.&șP��ܽg���%"o"ǅ���N�:|}6릑�(���Ɍ4�9 �v �X���B(�Fg�}�Z�I!�$�:�:���?,p���x��jh�+X�7S�Wk�+����*������bN�R炌�O�E�F�1�r-1|�G��|�i�#���n��i�`���=��uȇOu.��/S�%Td\91�접�@Ҋlʁ�Gx#�/�W��<]d�,!o �\�<q୹��k�Z�?᧭I���΍��[�w��Vi�M/����v����W����#���=)4R�|�D@W�o���8�^�sͺ����ΣU�/��g��<>����O^�R]��v���HI�<�z+��93]˚ �2�zMe�w�[��
�D$ۿ�恚g���d�ˡP��4?l�+�
�����0������9$�n��#�+����� ���?��}V#��� �b��W�)���"�ʔQ!��?LI��l�Z�Ӱ*<�%�Ά�� M�$�iW�h��Pa]�-\l�8Ӕz�s���0xi����6GЭ�_
�j�6�KD�������L;n�B#��1��9��$����Q��	�ƨ�:9�B*�'�U$�6י�J���l+b������C=���7
-MI�]��+��Z�Rs����ǉ�\��p���R��$ ��#���\zb�Vvp6|��.���niF��-7N�&<��H���O^NT�GZJԨ��^��Q��$���&4���3"������Q*�À�.�ڵ��}Š d�,aV���z����,��I��$�*`TK����F,��Ϡ�Q[�t��؀S�FK.�9���;�������v}��u� g����{�ض阯��'z��"�
���/@��l��|�~��U2};�G��4/����#�)*��+|�y�߈z���W�0�٫M�Q�-%��oP��: z���
�T�ژ�P�s���X�S�t�1���IP�X�U�4��6��<��hb�u�]UU3�*��y���)i���~�6�����6���ʍ6��L��W��f��4�Yŧ�mҐ�?]��VOGE�A�X���1D*,7fY͠ o�ds�?�����ݓ=6Zx5GN�4@��� �-��=��b'z��������@���!�;�a@�n�4�wd���	uXh�f�:��A�l|v��1đ?L%@�S��Ů�}��I5��	8g�:p�Ծ�N��.���|]�׸^(3�F���WKh���T�7�t[΅�s��m;Y�c!;j�������9<�X''��6K�3^r؄����?��o��8]�Q$O[l@@��$;a5j������v����E���|����Nw������:����s�W�]0?�V��%�&K�WV��z�!��>Oa>�d��5T3���ޠ��Y�N��Yy!+��g��8B�������p��$n�DZZ���Y��@���NļM~��8�j��t<TkWJk�=��n4��ֆ���?ӄ�/
+`���B�	0	Q�_T`"�0�Spأ���Af�[�*��!|�W	+�oū.H��u�)I��4��3�@p^G����)�r�<�9�!F���'�w]�;}�����lc�%v����;��'5X��9�n�o嵋�6���|ŧ�����	j�Zqo������Zi�vZ�5E���a�jDܾ�+�����C�/Z_u�9�]Α��U��wT�B�
[��Ny<�I�F�ˆx;���"�+CN��0�]���u�]-f�!�[hQh{��Cs�Y�
�s��^?�ӮO��v{6��#lݳl�07�a��c���@r	ӭh�������4B$�t� ^:�H��ix��P����{�Q{�YI���@��G(7�ߍi1�-O��9��FP��D�/���8��ѹ��?�tFR�������>I�=]u�/��:޾4Y1&��ح���Ԇ�F�:y��JN���~��lH�6�b��!帎ֱuɽ���r���TW����?���J&����`��g��W-�AO��mQ�Hkv^�4�CO������l��.��c�YV�CRD�5��Ϥ����2��W��^����DO��!��O�hq�Kΐ��(ʎK���ȭ*_�P�o?�W ��n�On�����n�&�wᓻ��l؛U�Ƶ2j�S(��1>��%^і�������t/>Փk��zχDM:5�*Nt nf#��<}:i@z`qYB��H�����:���s��)��zl�1EҮX^ �iߺ*����j�@=�*>�n�� ��%3ĴD����#d`{w�Bv8,!Dď�k论��9��ŗU�������[z,���P��"z���$}��4s�v`�F�:�heA�rmf8������Ab^ޖpl�Hj��{��]z��`:���#�LY��~�Qr^S&S��ت��M�2��7.��s�]��6e�{�r(�U���Q��?��C���bϞ����*nů��=;�١���Ȋ)"J�Q`�gg�� '�lc��z��^l��5�Cb�i��zen�m:ۡ��3���L��sI�A��"��+����{��6�B�|��;\.Gt�69�+Ii�m�S#{K����Z8��Tj�\���]P����L����mr���z�p[�N�T���G�V���e�x?fTa#����Bz��1��:q�V�]�nh��\r��BAY�v|[�\��a�zBZg��XAt�-�Ƈ��؄?/b���,��21�ǃ����ű�$1DI�nb��l��9�R��X��j< ~֖b��{�8��|^J�n�͠�=��h:�!�3���=��W	6�ǎb�1�l�����z���Q�1Z�� ��6>8ۻ���͸G�P�lc\i7�@����GUq�d�G�L���d[ٶ\�֓�+?�@JgB�x^�7��ʛ:��)T~`��:i�59�����X��@�y:�u|
��hlm��}�������V���c�!��>��M�F�.[�k�[�we���b:�̢�D��U�>�I���W���	�p�'}wx9l�W�k�ޑk���?�%b��	H`O��e*�B�&�j���Z��t�����"W0)2�@km^�Oa�Ag;�+$`�Ŏ���AY�;������Xd������H-��J%U�7���,J>��!8[>淾b
��sVO�����w������ȉ�q���TH���ȟ*�2�+����n2��,�39���5<��+��6�v����O��d�'��8�B�y�� d@��
/���ZT{�C����SB��aT����@-×�ifN��U,��DJ�[]�hC�9��k�D��f�Nr�����5?߀�Oau�:����	��� A't1ȑ�f��)p=}�:6�y�>�'C�I��@{�hY�N���ba�
�MH�-`*	��&��	�b�2n�*6��`0\-���#]���4tz�=OM,�P.�{6i�����)��Y��5E4���(1�I��5 y�<o�Xќv�p����թ�v�[��y"]��՜��s\.'���&�&�߬��'��*�FΓ<ݮ��3���K�=�1��B��zٹ�/�7.):���(�}�.(�V�ڞ���9��(E�R��9}.�f���eE�*������>�AKDm��cn�����}s�D_��k#"X�I�B�D{E��p�7A�*s�P��_w�6�3j���w�x�j"�>�����	�m�򣵉�p��L�_ԣ6�Q2���a�ܳuK�H��V��k��`��{z��3$
�Cp'�����;�$Ca��ܶɚ������pn�����"�aw���j(���$�x�8��o!�W���cijV��BI��'��Z[w
�f�O��K�O��RT}6R�+ʠ���Tr��"Df-�pql����õg�䠟�ct�f�ل��7�>� ���C;����m6>��0r�ٓ��6��RA�o��8ϕ��D�pq���t�Z���_�W{#����K���ߡR̪����%������z1#�_�n "��L�W�g���h=.݀�2_o	���Vң6���u#׽��n�Klr�]�L�ti�gvE�_��)&�VL�!��6DB�hi�n)�LBh��iUǮ���M��p���0�=�8�W�?Uu��-٨�&X�c6s	�1�-Mb��8ro7ޛ z}0�"�Ӭ�oS����lMK�X"���<`nx�7� ck�B��`˄�nIF�ҡ���Oӓ��E�(F��3�ޑj�z��i��2j]�d�M�s�܀��
;��P4_���ϱ�3l;�,��	<�e�.�#��;eJ7'�R��dl�*��'��K�c|�^=U�<�; �4�V�n�k*��Ǒd#�cǔ����B�@SX�H<��a3ɩ��6�[n�o!�3P3#֭����߷���TY�R�}�
���N�zy�EƝכ5�s�D.�C�t$Q^e�B߅�O����¼�Ќ�&i�j%�@Z��ޭ=}��D�}���3|����>.Y�X�+��F�N��/ѩ$(#A\�k���0�M�Y?w뛔nއ
´���^��`��)���>`����sS�h݅@����1&9͹ƒ�R+*|?�>�mv	�7�I�!�M6t"��=̖��a���oi�~�O���ʡ��u>�&����>wVP����.�6���A�xL�`0v
��I9����6U�?Ϻ���ġ����$,��φ�\}���8�#^v,j+��h�-ug��3�HmJ<��e��o�a(��:Hu�{f��?���Tm@h0//XG҃�=|B`��l���h��W�B�mI��9��
�ص^7c �@�\0~P>f���ʖ�#"�H�ߌ�����:	����t�Q��@���t'#.���h�DP"��暂�1��כ]4��VpYM.�̼�չ�� *��މ������l�8`W�DS�(���Ù]�{c�S�b��A��/�e�Y�c)XPҼ8%Z��)�y
UR6nD��6s���y��T��{ry�r�r�r�� EL�٘�����W��E���y���Z�r���8��7F�~��9��h�Nk�0{~�+�]�R���] �q�<��*f��:��9OG�Z��AmKq�Jq�Y-[�8�@m�Lv$�{�"�l�x�l�:5�Y�$���������~dh��"� B�$� J}ݔ�= ����x<��($켥t�$�;]]���],�ۍ%�Sb`v��5��յl�^�c��L=A��* w�?!���o{x�~6P]���b�Z�x�\7�696��xl�F�%����G�\~�i�A���n����3!PP����E���.���e( ���u���CN3��Y�D]@�f�v杖bL)l�f���ht�i1I����b�¾3q]� �\�<D���}n�tp��&����]��V�*<ݍ���8A0���>R�34�KH�
�r��1�G1����Af�����LGυX�!��8}��/��ib�~q��
����h���1�nw]@ ��0ŧ��tK�U���wK�ޙz�=���ܙ�G��}��o�i��UƤ�-3�n���:[kjڗ{6�w�}��|Gi�6A]c��-zzW*�[I�y+�����)V7�~�ڌ¦�I��O��4��<�fp���D���B*���,�o��6���=�gָ�& �����~L�^ǒ�e���c1ӷ��Fk�:�Eb+���?/Z���ׂ���#Y�eK�j���/�x3�A���e֬	/�U�������g�ڹ�_�ȺX�ퟷ{2F�aY'< �A<a�ٵBvی���q���%�*6Gq���`�'#�����@��+3=;r����hE�G��fm.���T��넭�ހ��^���>ٜ��sl���. ���>>����D�D8��-�3�,-�V�I�l��]��z�����6�=��ѽ/�O�e4����Y���@|��jڊb=v��	6��[��?j'&�i|@Iб��H�^�0�g�~~�u�7<��#��=J�J��P=�s������7�R��J�ҁ�,��y��BL�O;�@�ɱ:���|r�>�<VO[��$��oyGl
3`���}�G�����b�L��2�G�.�Ty�>fŝ��E�(ֺ���^C��D�{�����xb�(B?���A]�Xp�VV�/�+T�FQއ����zN��(��;��\�ީ�ƈ]��/��A32���n���š��{O�Y���-�O b6��>ϖ��Iu`4��Ip��s�(���ⷿDg�H�zm=��T�h�2�)����F���������%'::"��m��)��/Ԕ��k��"InR��Ue��i�F���4-�~)+G�q��a�ģ���E����OH�(����\�t����E�L(����7	��x�n�o��S�\V� �Gf<H�h1_ћ��p;ʫ<�[�.\H9=-F��;Z��A���v|��n_L��W4�;��é4��~�0�J���"Go��%=x��E�H��|ԩ��b���3N!�>z�{JMN�7m�ƌ4mJ�������`S�J��`������D��n%Ҳ���wl�X�Wb�'��&���D�L'��À����Ko�Ũ�y�=f�w]�xsN�i��G%��s@<ɬQr�1C^��>�F���-�u�1����-FKT�{�.�|d�'���Q#&� 29#�>NM{��s�!N�a:�<c�ۜ3v��Tۺv���tQP���X���?��(�j�Pc�8z��(y��r��	���2f5�����Z���t�c����nSh0ߏk(���,����v@�y!����g)?��,RK���ТDQfL#N~����YK9�Y1vdv�ۣ�q;�w��5�$��ޣ�Q�=	=:vb����V�� "��l4��6�Y|��xSU4�w�%<r�L>?�M��6u�� "�~[Ů�H�t���~ ;�r5橃7���q�ѓ~��t�ڐ�Ld� �+���,�l�X�*:!��CQ<dz�]w~=b4/J\J��p��-x�����3�sf7�j��m��@�4�;iM`@�ͱ:� !�5���dG�[9��}��]D�~��2���D�P�0���2c%.�%����e�n�'���# ��g��L���<r^gÐ��C��]ǼE)E0x��D�ODaë�}��=y�m5})�}$�pb3�_孆,��s������3t J�8�d�EOEG�HR���Mr�����rsz��A�w�]<�������U���kF��E�� d��"&6��%#aN:u����|�	������VN�	,�*�F�Sb�ȁ�,_W��
�V�QC�*��b��Ԭ�ArT��hY �����Kk&yҍ偫w*	4����|x�P�E��lu	� �ُƣU�W�7�R�Υw�.;YiIrJg��0d�4Pۈ�3���uZ��
Sa�Q�E?i��s#A��>Ғ��T��)�b��Ƌ����&�o=��U���1��0R8:6�K���2�+�u��#Ylr�n���~)?.q�׈���M�'�w��e���K9GMi+�=����i-Fa_���}!3�q�f�'��v�����!�0*�DغvX�ȗ?!D� {*OjY��L���I^�[T`P?�f,�(�hUҌ�[�")�,7�*��iJ�^4���k\瘺e��.��#'��2�I��\}_3>JV���vF�J<�z�c��؃[�[��S�����l��+���V��X����@y?M�7B88�C.W!�.]��mu����)�'�����?���;7��݈�\�F��W��r��� ����'��'����͋q&�&yC���TI�H�{I���zmG�Z�vG�����$л���� ��[mI�W��{�$3�Fj �Z��Q�._UE$Sy�@��I�9�k,3�"n��H_��՗$�]y�#��k��O���W ��`ɶ��ߥB7� 8�Z�?�zJ�Sٟ{���E}��hh����&����1�*{�}�)��]]R�Sm#?����%cIr����ǳ�R9V� 5��'���w���1��&�t�jҕL�|R��*Nql�<�o���8���@."G�'���ϧC�t��-�ql4tR�U�n$]2�U��W�آ���Zy��<B%�3x�.�;F1��j�}��<��彿�� 77���}ߒ&�����kN��bc��k�q��D����}^�W� F��L�,-��b`E�۴ר���dk��3DKA>tgo������|��̨|A��H��y�vsۦ�s��-<sL��r�~�ȫ���]������ ǳ>�B!��h�� F������DAnt�A�r��gYY���F����v�Q]0.�
�ȩ�[��C�]
�]�91�`�e\�-���*��KKה^�����"	~�tؐ���؂S�F�.�T�8���������Aw��z�?�	�X��K��i�w+m:���]m�G���P��� ŉ� ڪW�Y�E�����X����x<b���9z��m�o�VwyqS-�I�e��w�65£�S/׼���)��=�#�k0���>J�ڜ���<!Z2^�[�z��P7�]h��Øo�,���/t�u_n��c�W�[>Վ���%4�;8%ʒ�J7{|CR����N����_a�.&*�+�hZP_�h�Ć� �4]D�L�L��$���銷߉��ĵo�����0�F����ߜ�3�£�������J�YL� 10�(( 	_��x�%|M1FV�)�'�{�	Ą���N�������St7J0�.'e��C{Wi��jj'B�j?��	���:���0}a�v���n���a�^0�?īd\B��^���/sZ�I��܏�`�
�u�FRfb�+�w�I͍���8��n޶�|<��!���.u7����RM�w�@bM�E<�{"�*
6�g� ���Rm���1K���1�:�P ]8�c�$W)n�q�:#"3(fނ^W��������]�.`�&�����!ov���r[����B��v�Grwi3�1�nP,	�~eQ�����ƣ�S!�ѓ�I��D_/�W;QU��i���6�8��}�դB��I��3/���ĵn^A���T�޼�bc
���]�o��f�V�3�>>���6rH�>���9k�I��)ch���T6�p��[X/g�J�"��!N�h��!���h�v� in*�q�22 ��]��5(�!W��.c+���Q��#28X���ŹDڢ��(aoߙ�EΙM�?���[ӗ�)���7���m���S*�o�"8�7yS��#3�u��K�9$�Nc�Qu�X�\�펱^s�Gk���5^�?Q��R_=�aHy�oD4��w��}'B!�"#rs
�ἇ*.������j�+h5���ۦ��MDGog(p���^����]�I������������YG�I�@��Ï�Vq�ICi�m��=��Y�H�^�.�"Rˇ⹞Ԓy� a8�_)�S#�����Uݡ.V��A�w�L@J�=��ɚ^�~^J�_P�	���l�'�{j��l!��w�U=�%�S�l�u�����1p��1U��!���Z3��V�O�$z4~َ�ɑa��25��=��5Oh(��K˷��^���X9T�J�+dރG.^�~�'"�g�ɀ�k� �h�*>?�%�N�S�g~�մi��ʤ�Ƒ�]N�S���P3aRv�z(3��m����U�o~�;�&�RR!�W�&b���3�Q��.�N�3ڊ#=�6�6���C �1eA�Z�K�&:8�	����:g����������/W�(�����fީ�k�Q��V�3�v�Ov���X�I��-J ��Z�^Rq������|i'l��l�rgP���S��p�(d�I�陭��i����\��8*����'/�)4n�0g�G�`���(P�ȀJ>�"����1�0ڪ02���rL�56�Aä��.ۏY~S���-;��f���¹�)M�<1��P<>�V F�Z�:���U�F9�1��l�ŧUUD�xT��j���d��]z�F|N��+�P��?D?�u�L�'ɫ�(���7�)���h�2�O�Ԗ�cׂ^$T�Q�_<(+��us���uQ��@+���J'�Z��C;\��ד�yV�#��4FEKPc�(�^��?�h4������@��.��[�ipZX6����'��)�Qf���Y��|7��`�S���	sX"�E`��s���CN��+L6@7[����W7Z�0fy�#��=h�% :�	��"�L-(E)�,E�:���PC�3�y����2�
w�t�/k.��ﺍ,�	�zm�����t���0V�g��	��}��D6�/��q`ę�p��y��yG�C���"�v�<u�#'��z.�~nt�!fw���@(U�N5�p���G(I��L;CA��
%wJ�G�#ʢ]P"Ε[����I�'5���ᖚ���L�
h����G房 ��g�R���$��3-'*�I��⭾�n�P��D��׭���pI��se���v�<3Wu�M 9�?����E2��@�h��x+�J�c���1�V	��������[v��:c%��x�A����o�o��p~�K�gТ�sj�2��G��sSW*���mz��/�;:+������X�<n��PB��o(��5�������o�>^{�����	Z��W�¤��𷑵�:	�!1����)=~/�P�c��<,ʣI̬k����d� ωT�p�Q�u�Ų�M�GVZ�Σ���7B${�	��;j}3UI�IQ��OV��Wv�xd��1�T�2�ex �ؼ��\���(��W���2����ln�=T�����g�"�Y-ҝ�?��K�_d�U�YqK�G�~S\|-�摲 � ������l��$Z���������§E��+<�����@a��j��e>!�߯����x��4T6g��
�9K�1�9 ��")Zz)`�1?����סZ�`<a�|�d[��[�YT�6�M��l���JQUz����=��](*������8����XI��F�� �s(<=���M3�`�UA�j#>�B�8kT8�	�%�7?�\(}pČE!}�
 TZ`�*���Ҫ�I)��Iع��%�b4�Va��L�mŹ ,<ޞ�sm�
�E��$��\4��Y<�j*��:>��� ������
�j��@�{��h*Pl�<%��E֞�r�9G	wK3Kȝ�b��:�����<��W0�V�TG�h���7���Eݫ�=FNw��r���'��NH�������?�:~�����A�G�֮�| ����tYɐ�k�q�
�V��%V`m�a-h�ґ���b���2���R4k�t���SY��S#�7�t#4���\�5�p�A�q�N���R�Et��p�^�V�s�j��nv����A"\�1j(��-*!�Q��>}Df�а��ϣ4o�nVy�@�e�m6t�-;�][N���	�Z����l��>� �aTp�_/��o�^��nS��;��/��K��D҂f��c�
*����e�L6��
�9�y�V:-�Qy�)�]G��g�����*T��D�6����ٗ���= �	`Y�d�*l�R�K&�9ѡ�-V�T����D'����ẍɽ9�jJ��@z�Q��I���R�x��\�D:=�X$:� ok�~���7��±�[���lm(A�����ݭp�#��`*diu��#�re�jA7'憇��i��ڀa�6�1W�V���fW�{$I�>fcni�3�vȝ�0��tQ�/pccxli����)y��Cc���ԏ"�)9��>bЅ��|u���;c6�_]B����m�#(�V�L��.�#%��3�0��<@�{Ӎ%���,���R���#���Ҟ8�g߬�'�ɲ 5��&���Ӹ��ً����Q��%�B7�i��������NMU(5�Mmµ�-�oM�-c$	��	Uo�\�W�bܖ����~��+���
��y-Y�s�!+�UҖ]�h�ùO�܊��P3l���W�ҭ��̳���X3h;nr�3��N�U���il���o�5}�f��?��?y���p�#0�4o�kzͦ/�=?2N�@��VC�� !ݚX��l��T(��s�e`x�[/�6T�7�)�ƛ��8x4�q�����~����ST�����G�u�߹EU�v�+�C�v$A�!�,bT	��r�\?�̓�L��p�l}��!?z��g&�L�W���0�'�9�^-V�ܫ�}��酽�~��&����^ S.:�BA���2���X=�����8���ԃ"�8����@���������=���(1�$d� �G���k:��Z������C�f ��D��\�YU���ť0�9�һ��;\��G�a߅9���{���\�U �c� �	gT�ZIl���4G���IIw��`��,;�kJ҈���7�Fg�^J\C��(l�����-]ͬE ��	���P��]T�Ũ����݅�E^��:���Ki٩��S�M�b�$��rg�t�\{���E[I+����I�O衽��yNl��LL�9��NF�������@�]XQ����^_�G�Ww�yumܫ�ڏt	x33�����UT �|G���ﯟ�t�����-4u���^2!�|F]%�I�\k<�v*rD���}�`�.W���wV66Ӫ�Z0��l8hA��>`��b��l�ě�Y�e&_+��G���e�i1���<��v��Z���Z8�`mYԐ�e�˅�4���ai���\qO�N֙
��|p��m(fo����4<Sn�.3��T�Y�u��5�dy�I�8ۥ���L2�J��Z������|^䯼�,ȷ��<�1�6POmmF
����.���>�M�#�ͥT~~�D���lgL�]yNiz��c�-�����z�E]�E�=2�����`�C�n�|��P��nEY�����\ʄ�Z�Go��q(�}�N�	�8ܔ]b=�}��G��S�8�,�k�WHv�_���ï��99��^GFX�N���@A�@&TKc������BV��yȓC�}�V��L/�7`q�ҿ�a��������Fى�f���7bᅏ���ʩ�P�K�2��9�z���d���]����^��"T���f�k(��x�=������D�E����8~|��}�4R�U����v|�������m>�$��	�<�,r��\�C�,K8г����vœ�F��N�'pILQ+���l�ٗR�_��Ӹ�#�˓��6���l��
�r�\�˸��Y>֝�O��C3�t�8�q���Q`@�ɗ����s����Raw��n���e%[�,(�rP���&S�c6���yN�;A�'&�Oe<s�S�yY��;�`��Aε�AJ�)S�v%ɞ8��>��ai�y�z�,v�3�PGU�A�v�1R�i'Oh�Q3rD���c���/�~�!�0���A�(̟���k�����ữ��:w[�".�@�1��sv���D'����p�߰�껶�#�9jp�<��#�a��V#��Og��6�w81(�(�܌�snq7}_	�N���7�"�Jr�N�I���W�V�����{�y?Z#��3�ېF�Q3��k��I���Ў�핺�h��N��lasyUe�c����{��B�Fx0��x�>_�}q�RU�x�T�x�މo������sk2�įL�'1�kzQ�T�ݑ�J^��9�jT����B�*�o;�N�zP�ɼ������²�z~��dT�+K�'&6��u��zl�F�����)z��i2�q�\�s���m�S��Շ	q�в�஗��:ٽ��zh�j���:��Š��}b���J�U0mF1����3j�q�b-�>�/0�G���~��_5`"��}�O��1DbY���C�&2)2i��R�*%׍���@�}e�3�(�ݥ*:P�5��Ėi
ī|`J?:����l�tո��8�F��$�8���` P�����-�ht�槞p\�=e,Of�Y�����(�ɳ흃���)+� j���'�[�l\����=�t��f(j*[�SPn욭s���_�;�a�RfSD��5r-���s��V�,Y��%_H�n�%/�P=m������핢�?J������g&�8��D/��1���T�ʘD���-��(�[i���w\&����5|�!DVj�;��%��X�������f���hLM�-�\E?��_L������]���2�����g� YK���&+y	ÛiDy��Uu^#K�����g��{`�VH�R��w�����$K���a�r�
�ouSZ��p/f~D�%����cGѡ���t�yj�=0508��I�D�7��"�&�z|�竈���JЌ���6~H,��n����Q�A�|���6A��USn7�26=���x��!��R�~w45+�#î�ύܥ���p��^�Ğ{���{`p��Z� ��M���;����n7�7>?`>I�)�+V.��Xa.��x����~�8ǩ҇�h�t�c�/��9q���eb���:8"=P ��[�
�ZxtZ�O�V��=��B�/A�L�Bz'���4�`�$�uR{>�D�';�s����\�5jJirx���mub;���:2Mt1d�wy����᎗#�4'����[�&�]|�r3U���藳B��j�-��Gxn���r���O��Ӛ�K���=9п0JH��������,��+�����;r���=G"d�ag`�j����<0�(��c|c^����� sȅ\ʲ����n�4�ydض�	�7��2��ߺKKz�8���
",M)�ɸ4�#���J�U-J3y�pz�L���]�.{�ba��^*�L3Ɨ</�(g��^xob!X��aI�_�3(6	����4�"���DzN��Q6�lw�'OE^Z=��n�S�' �B9Gp�C��u�YM�দ'6�D�f幂ap�q���a�2�ē?��#��	�6_��p���+4�$)�Y�Z� �;�v��9������p�I��w�+��A4���h2;��u�Gm�j-ɖ#�����������U���X�'�h�cAZ���R�|�E	��E ��.=g������")����p���\�����Zn�{Ϥ�Q9'� �������M����x�*ݩ������sf���U,J�]�c�P��h��'�6��z>s�i�aV�:��~&U_��4�}�t@���Ƿ`P�4u��/8k�N�
&x�5����o� w� ��.3kY�����m����y���1�c]�κ�]K�m�����E�2��++�JG仅�����`�aA��4L���Bx\�)'�z��㴁G���)#��ds|]Zȭ�}�W����+0�R$���&cY�����B�Ȏӫwߐ����\D��ut�O��%!у�=��z���c�Ҡhc{�O#���9M�nT�� ~>����� ~Lv&�D��4��\ H*�\3&�݇��
�d�3ޓW�Ii������R�?�f�7�'�`�`Î3(9��?[1	[6rC!/�kd�{���`}�]����9����a㆞ u�tx�{Pl��J��2���8�-�M%�naۧ��|���Э�YL���<b�����K�V��9���AZS���E�Nˬ���Z��R��&�$g2C!���@�[�ڨ��g���]p���v�t!��]�_����7�����xF�XS��#!�k��� �·ҵ]��^��ޜ��>��7M#:��P!ezD�wj�Yi�}$�~P-��/{���_��rЧ��������N��Is��{�}{��ę�U�N����Mk䵌��� �PX~���!*J��C�de�ᝪZ����^�/�|�Bݪ
��bo� ���dB�6���|���mj�<�i�U6]e�.�>Z��UP�0([-\Ѽ(C;�[W��;w@ �L�� ��Q'j�Zw%\9�ML+,v�+^N ���瞔��u	Eͽ��!����!-�F��3�(��%�-��,�_2=ly�fs�f[kB̔k���m��!�--��̀�j���Zh��f	��y�7�� ��HC���DɃ��T.V���� ���)�o�2��B ��rFԊJ���]���F淩�Q
�)���b�|.�*_ ��_G����P�)Ì4���(Ϧ�\ ���))YWV�^�xB�F���7���y�� =#ufgQ����A#9��x;/���2a��h�nV�T�w��ֳ��G����$�'�^����Q�*�x�E6�1�>\R�C�&��84A(��E���<NQ^�ޓ1(�W�z������L��&�
"�Km�;���C?�%2���Px�]ż�xnp&��ڑ�!B�\�ػ���Ț���gLRu��#�R��8v2�1���~�_�Y��8�Ī)�������
� %��i��w'q����k��y��_��;V�z�����:2�(��8�k*�8iQ��;�2������hZ�*8�+i�Q�����A���Y�� Pw�
�]��=�VK���i�=�fP��\�!;��'�JT7^�q��U�"W+��Y�M(���j�zNx���x������_���ľ������)���Y�;�?�y�Wr$'��yx:[�p1��F��̺��ǕYuC����'k�l�*%��C� -۶�j#V��j]ltD�tc��-�g5�?���`�.��2N��|��=����j�)z��H7GI��)��sJ{�xQ$�ȑ�J �'z�./[Š0x �1Yv�D�e�nّ��-Uն���M�zL�o�H]#BfyQ���^��IT�W��$d��Z3�$�l$��:�
��3~��ů�T��uU*\���छ�b�����oe:��s��N&�z��L](�/��ش/�/�G����n�����~�=���_��M�� -ͻ�'����hrq(/���*Ũ�N�����ѵ����H����9/Z]c-�-#E��`hf*�e�Hh��䞦��Q��tC�$����<��E�`��r�3�g�h�\������O���m��I>t�u��k�F�'��(�
��Q �7�4o�u&j}<�~`W����9�ƕ ���G�>&lI��{���B�X�w����J��GTǦ��#Ô�H����W�l`�W
(;ߒ��j&;_'K��8�m��D�8���C�9 ��),
9	FO������}��&a��!�x9lYl���\E����+wĠ\�xm{��s��2r�?����D(���5�ص�N+�=�^� ��:dK�9:��m�Y�5a�q�R8��4�{9��#�@��6t�@�kW��r%SO�ѾH�Z����y_��T�aW�^���(G��	���Z���0U�, �o�}�s L��r# <��~H�ka��v��}[�!͉�?��R��m�ZH��	�;f?����*-ؙ$|�����Ћ��h�����J����$�[ͣ�p���v�  �j�S��j;c�s O츳���k#�����݃O��V����'��M�x�#�7F��ïF��`�]O<}�1}y��q ���fs72ݽ���
:ǅ����f��(�U&�J  ��85xe��1��{�2�\��^u��P�ɿ��O`�冸:�w�F)�4-%�F�NB3�h� A��I�)�.k�F����G�Vp�F�w��`Hp?k�̛ɡ��[F>�s�\j[��c���5�j�Ms�q�u�2OG$�r��}*�Q�S6�[����N{�+ ��{&�.�X�/��}��R��X×<�X$�Ǹ����a2N :^9���F�����忩�����yJo����������Ӊn�/�?R��]L~�F`�/�#�$�@��=o)���W��J�K�N�+�U����(��:����������;�d��q��:9Pǿ���Z�@�H�%�w�D#�9t��M���#��%�J��n��5���x�O��� �{HwxU'g�*%��bmC��E���o�j�o�fy(������z��t����?ȏ�U��j��x�ϣ������X�0~�4�VC;=�� ��CaЬ�'�F��K�������trs@���J}�Z��?��"��/�=�y�f8ۣ�Kij8���uY���*�|�;��W��!��J�N��b�7��3>�#60b���6{��Z"��[�>�E�6T�,ĕM�+�����NaB��H��<y�[�^���6Q�;�"�L�p�MѸ]��fY6���e�K�گ*{Q���y!_]F��T�X��%��m܉j��O��gK_K�;���N���l�c��������D��y�nR�	 r�m��P@�]�ֈ�9sh)��	��!��BE��* ��	L�F-�Ʌ�r�<�I�:v�d�[�Z�W�yM��0�!+iȸ� 	*D���8� �O��*������A�Ű�kǳ�w���x�[�&���;X�Q}Bӡ��35�\�xf���Kx-������$��|W�@t|'x��	���Ϙ��E�`��>��v����nQ��&)I��׻t���U����w�������ov��"P/�!} ��?��˚˝&
e��k�\ҁ`{���ٱ{d�����Xm�Wϑ��e�-�ꏘ�ѣ��_/����n�I�8_�)#�?JnJm�}�����l�
���j��N�͉T��c�oʣ���B�lm$�8&lR͐�.���AG@���c�Qe�]�p��CYɉ��X�-�@ޞ�4-^���VciDv�&Zy?��l���v؜ѿ�(�0����0� ��No�Js,�@hA��L6��0���d�@��	/kN��BT��T��R���[e ��ŷWL���TXJWG?�����V7
a��}O��U"��Zߗ����҉g����a+D��|�h�|T؏93|����A�,O� `h�U��X�T���b�iN�$#�Du'�h�/�/=��CjS�!'B����qC͜�����C�o��i��>���f� u'm�S��Շ��������`6J���jnᖋCJ��X�2L��cGՌ:���G.I�Xam;�d�����.�DH�e�h��o�PyH1��>�Y+����r�D��i��2g���}4ˁ�&Ő���< 7��0�~B�j�y���##�2���@=��}�J�c� y�'Xt���q��y�6�>󞌰�����0�ڥ4)p��rMn���g��>���ֻ8���d(oQ`�N4�	4)T�|0x�:��S��#�������y��KǇ��NŢ�T`_6_I(�k��`�Q8c�F���ɔ�珔	F�/?R����^����X�2���Z3��=?�I�xD�8����k�0��)�r���R�%8rǏ\��������Q��73-����3E��0!�˅j��žW����O:�r�;���mC#�� ��{��������y:��SR��k[���}	�;I��y��&���;d�����d|��ש�	~��Lg����hL���T�30d�l(� !�Ւ��Dn���]���?����PKL���#��+��:YtV�i�O�YB���(�Ձv/�*�`���fW���D���+~G��7d;������r���GS�i7�?h$�t���yI�R|E� �v cZ#��78���|�Cԋ�/%�kd�͛�����@W�Օ`��>�N���j�m!V(}�6�>��o]3�ae� �*�2!{���)�����&���3��y�܅l<e$�������+3�a��g��F��T݂lDv���H�ÊZ�z��B������oH���"�¿V����D���B������(��?Kh:RbQ�K�HxJ�������w\8dtZ���U���!��gJ�������Dj�"����p��h��	�6G��{�n&90��|�^=�:�2L�͇.[O�Ę(��v���T
���*C�d���3V�;١"�=:��w~֒�7�[���?���	e &8!Vd�#�f�L;�hH�M�:�� \��������h;o1��)e(��a��$T��>����3kD�UA�9�J�Lk������H*��*��D���o�y��>�:�w�Y�`��ǡ��A�Q�	���^P��:���,�з+��՟��L�0jz�5�UN<������gN�:�x�>�X3�'4�#ڮ�{/F�\z0�^`G�	������-�#XB-ich%ϱ�PW:,�b�-{y�[����-���qe�Bv���{�[�ʒZ�24]j�����s.i&�<mhx��C��A�H}�8Z|���˾�i"R�t�pA���xE��ݣ�.�D&O]��jC.�ks�q:�1���u|���Ui9��.�R|tt{  �<���C�e�{:j�%k<'~<�;OoQ�=d	{][�~,�Tk�����-y΢�U�!�AI�,����1J6G��Ä[�8"�AJD+X�������x/fتX�\���Zw
/��{0����Ӂ�T��wLa��u�ً�x�7ܵ�\�g�5�݄]1d�'u��L�~4'v�R1G�Z���]� �"4��l>��g7W|��T.��%��0pI0��"���TƟ�QJ%8��/�t�|�k�6_.�f�����c�'�~�y(�7�1¢A��J ��Q����6�IhcQы�n�zS����;��[͙ ԯ@8d9M��4GpN?���)O��_/~��	���h(�g�6��|T H������~�?���~�`6�5�w�Xl94�aK���*�S�D��a��K�'�s����[gT��:x·U��1�:�Tl�Цu��p��ScN�{f���M���-t��~����p�vBz�p2z�Gąϭd�,�@�^�	�:��e:

�X�)�|;d�0���2Is*uI;kU�5I̅"ڨ(,v���504������+�&U��Z�0�h�K�ɇ�q�@/�Y]�n���};�AabԼ�~��ba%����,U3mj-����+�h��D:Ó�M���ߘ`�N{���Յ�#䍠uM�z��SI�?�]�^��j+���aor��:��k�Pm�`�u�XPi�q���R��3���o���Uĝ��{ �����S/nBM
�Q�|X�`߾)=-��e��rr���q�4.�J�
X8���nO֧��F�����S���
�� sS`�X�1��C�W02�I8�c��H-������(�`�Y��VV�I
�g�|%t�}\��/U
���3��Ǆ٨�֓��8�" �n
KI�!ʗ��g��=����덉�\{Y2
&ϼ6X<e㏥�M!-&@_p-���O�����A�8�w��~)![��	Ŵ�����Τ6g\}X��`��6'�̃���=��/0��`����Q�h�	�K'>�}��GRw�z"�u�X$̑�xh���_߆DpRch-�ܓ����Q�Z���dy���]�ޜ��Y!�X|�On
�3v)'�QZ6��������H�>�_��ċ��,�U&� �&<����7lP+���$���1a�)!y�e����!�����"�{��ۇ��u~V)������YΡ���掉���t��/���9^S�Ap��f�:1��,��:����JI������U7p������7k}�A�o�Ȧ���c���Y���N�R�_�����l��ޞg�����9�P��+��cQ���4H1 	}�jF��&��J��*��,�ׇ�-k^���ݳ���"=��"X�ߺ\�j����_�����<}�!&��8�ޯI�0����F]q	V��fZČ�%AtZ?��������4J,CQ�w�L����8O>_�p��:�(7���TL�>q��(�F�1�n�J�(��gs���C��*`�z6���q�\��Kk� �N;�b��^����a	�qvy�~�t�'	
��U�B�p����UDy��q���]��]�rG"3�)j��C21�cw�}�)��,-��^��������4H��^��=B�Z�Z�C�T9��
D�Ys�Zn�5# Y_B�i$hT=ܾ�8�;S� �T�[�4+Y2�Sir�(\�ʰe�<�T7�/���+����6'D�a��ۼN�{ne�I��㼗�*ϜA���:ܐ�}�E���2�]���Dٴ�H֏�L��@�H�_pd0FW����K{�������W$)ሶ9����x�x����[0L��W�n~UKƮ��kt-b�Fw&;�}IG�cGP��6a]u���f�[�FW� �i��_J]=�	�p�W(����nJ�^�΅I�*N�ʉO+��s.N���<�#Ak�vP	�Xj��~���i 6�R��m�lQ`��ƃN�h�dt�{zT׸�aʫ54��{�`S�M"}�7�oEe?��1p�3.cGˎ�q@�	|��7l')^�#�N�g�65A�wx˖Z�٧��^�~7 u�c��R� ╊����_��;���N�!IB���N��F�@�G7�9K@)�*���믂"�C���x���B�Z�p���R2����� �"��fg� ؙn��Փ�j�ބ~KC�<S3�p?�$��7|����q����O�S�_�2����x��M�j�/ԡHi��$��dȺ^�� ���.@O����j��KӃ��;��	�{�e	���Z�A�d�𮮌9	�bP ��c׌p�T��ߊ_x�H3�O��|m$Q�s7WBe=6��U��9��.�uD���?�8`k	yx�8e���g2-cU��`'z⽟���eӫ@'��>��dx��~�{N��1�������8���7���a�F�ɋ�0�3���j e�ё�Jf5g�y@��ծ�
DGN�\x;�nաơ`V��V	Q����7�dR�!D�(�S������:m�D�7T�c
g��U��A
��fn��z����4=���az��]���(�^�c�q��}��$�흸�6����7�y(�����8%�ɢ��y��T�ϖ�|��bA%N˳a��[P�\�zi��M{�)^T�P6!f��e�ꎼ��W����������|鲻�ʤ��6*.�����#D��Kػ��{��t�z���n��i���W1Q��8�����o�:j�N�  ��.�P�n�	#��Fǀ��#�6#������ uhp��ɒ.��g{���vu��3!��\?@�?5`�g ꮾ�����Ҙ�5\�(B�g�� ޴~gp��kG�����2qZx�u�#�~9�|���V���c��7�͠ç��\��?�Qp{�4ɞ
v��t&�<��N�����%�
� ����U/p��������I� Rv�aYq��Z�BT�W���3Yޔ��k�ي|��I�Ǩ���
l�ӟ�Pgx��P뀬)��ԍ��Q*B@��w��\��葇Rh�N�Q������h<�0\�3�di�4d��3l���d�J�-� ��1߈��r�1^����˨cm�r�(��9_D�	I;LJ�.Nߦ��}֑��i�꧶+�*�9� ��jD9�F�5ۼ� \禔�-�Ӹ�P��������B�p(�e{��\]U;3�W+�u�e�ܞ�U�]5�U.r}�f���@.� �����i�8�^x�sq��\����?���PB��f�Z�!��1�4���@��2 �Iri�tp��z�0�� �B�����e��LӶ�����E����u��_��բ`5��;c�u��;�ߺ�r{V&�|Otc�݇l���n<��fhTm��)u�[�BV�+V*�%`����
����� �Л`��$r3�`
A�sF��ը�2�G܌�WM_<��KX3�^�m�r�����&�8��\�����R𫔵�a�g�2�V��tx�JÛ��`~���"����u)y���p��'`2�{7�G�+К3��� $��t�"�����mHs#���M�O�.?QmzE?+���d[�3��؁9�0٠�����e'�of��YoKɵ�-'b�+_�kk��He�f��9��o���-0��Z�m�資��Gm��aZ��}'n�n�֫�`��q����9��ʵ�?�����`Wאԃ4\]�hd�L���w��>���e$��^C�/��r���/[��:?�R�o���Y��׉�jt � ���.qv'�A��b\Z�z�����᫘h{:��h"4tAW��Rj:�}x��Gs��7cx�!@�z�[	Y��i�y��Ѭv],�X�.�(L�r��H���ݞZ(��r��Q�C����y.-,�b�5�&�T���^$�R,�3�dĀ7�`�6��Q@L�W�ޛ��$��IKɦ�������m98z��D��SE��|#1�k�(��Ă0�{k�2������u�+�H�c5������7/~�9�|}F���Fn���ܾؿ�0ɵ�
h���K(/|�D|�k%}h���c<Z94rf�4��H[y��y�$V�S����(MQ�f?�����-�W#t�P�; "-]h���֜/��mJb��y$�spz�-� �H�^t��A���4�v�{�ޢ\�g�������>"�C�s�G�Ơ	�<�ip��|��*o�b�B\���B/��������)F�T�M��]}�b%��c�PU1R���#� 1Ć3����f�q���,s{��eZ������k�<+L����y$ߟe��5���C!�%w�^**�u]q�S�IB<t�I���[NbƅC�g��:��e%�\?<{��1p��o�t6��v�M��E�k�t�{Ֆj��Z�`�1Ԏ��?������ޏ@w�YR�l��805x]ș�?)�<����{S���#g�9�ؗt�����Q�4��z�	��<%r�����E���i1/'��cR*�!3Hb^+����e=����F����^�f���u]Zs����>ϱb��/��Y�o$x@D�%s0{Њ������[���f�g�{X�]@�1�
�^sk�RV	�kV�x.үIl�@��*˳ѥ�qym	���"QlZm0����4	&�i`��s�9��xM�jp̪5P�1R}1Vcq5Q�O<}8�v�r!*7��kI"��EZ�,���� ,�9����e"�.j��-C�)U��1��6JWK����^!KD�8�V��1���]��7� ��mP�~��t<���}D�F~�Q����y�[��$`�<�Nw3��ݡ[�{6��b��jeI.�����$��hƵ.����TS����pe�0�e����${�Vu�e1+�P\��%��fܮ0�!�n2�OTtߚF�ѣ�-�7O��Sya�Vz'���c5�Q�(ګmxT�J��U��_��A8�H���3��I��%|���ܤ��ϣg$*�翯�'���%�X��(�"W��Q�Y�*$�c ��!��fؠ?��>v��ѥ>��Q
�c-�2�ڟV��EE����-c�MD��D��bm�����}�ϡ=��5����`E$��+Uڱ���|� ���bI��SF�_e2��?E7==g����-{��E7�m[�cc��i��uߗ�x���z]�zjT���44c=�z�0.�x��t6Rͨ�K���;�!�֛���Aӕ�p!j3��!�{ĝL����遄�.��Ⱦ�_�}hB�(�V�4��W�%���a8VƝKD��l�τ�dɤ9����n���NЁ�('�!�'�YB}ŨY�.�ad�����|��mO��ґ�2Ĕ���Ŧ�-��@C�	��i�ɓ��z'r��惈_�a�����ڑ����G��r���͌r�Y=rnx��D��]m���G�V�f�[z���7%���>vi�u)P1��p��z�ekI������V31,��_��hͦ	����lhzND��o�o�/q���(�_V
�ĸt.cv<�`F{;����usO�A?ù%NjQ'�cWͤ/���m��j�= �'��<�35���.��Ł+_'%e�"#e��W@u`�^QJ�Фs�)TZ��័�Z;b�n�k�()m��%��4T%�}bB��
�I�|��q1%�˨
��LN�Y����F�*����SO��xZ�	�6A�&k���L>�tѵ ���[x�� ��{׽j��կʇ���
��UC��������A�:���L��!7ס���@ٺ)%dZ��e�h8Kc����,�ЧS^�ntk�;�Ѭ�����#
�1���A�Qh>�]��ѐ� S&ɖzD7 ��ӇO��C}.�!|���Y�7��>�3��ya��ރ�B�d�g�/"���x,ɸH�S2{�1�bӸQ>v��MA�v#��I���su�����u��tl�g*<�O���gd�c߸)p��wԑ�5M��2 ���\�һv�nD��f�wOڎ����G)�f��X�'��ʙԤ\�\b'"�,��p�c�Luu⇊@�I���4�����'�a�?�`����NB�9���߆��Y+��&��܎3oM��p�z���ڽey�MK-J���0��G�,�ŗ�#��㢘c$�~��K�̹�-o,i#>+�M+�o�|�����o���A~�L�k�0�wi�=)���b
�H��l�Ԫ@�%m��䭳�\.l�
�i���e��|��p����w�R�i≙Ma�	����S���R�� OX��~ǰ�%T��[�q�H\w���ZFVW��u�M��~7���{�f' +�F�y���o\ V"�P,����F�8L�?�H�H�`6�͎���l���˵�1���B~�Ҭ �c!�)m�aOm�tqJ'+N��T�E����Ѭ���n/����S��F�5}d�ckUDB�d����|B�c\��A�[]�.?`�7�o8���`&-�EZ� ���?=��g��o/ �p�|���m�h�W�ɺ7ꂁ�[���$���G۲Ԙ� L!�����+�૏>�q4V�D�/��g�2N'H~��%�i��X�#�ĤrR�S�[�.4C=�N�9��Ԍ쒩EоM�z>l���f��Y:����@·-����8N�ƍS�wN~U��e��\�`�Z�wI�*	v��ݑ=�N�r�Ew���� ER7�6���. G7���|i
#Q�����;�"Y��ҟ8�d�4F��f_��>�W�;')V�~�Qv�?r�R�Q�^)�]����=��ـ�P��٫uf=d�l"��v�?�D�c�R�Ko��F$z��ߛ���J��N$�&!�ѐ�����&������5@��c��?e��S���w<FQJf}��ճ�O����]�͎U�!L��Z#s٘Y�N������{VCm*���v��?|B"i�Cy�
5��T��p�V:�9ͩ虏��'Y7�%�έ�g�vҠ�w���~����#F�B�GK�
9ȵ�j,L�&��G�)|V_l������dL?�=��8�ܬT�U㘡˥��$o��-UKU�����8���Ȅ �V�pщ������u�i������ZZ�M1w�0<6�c@y���s!]#��Z/X��^c�G����eQ,��Q�PhRg�s�IFo	!�g��8ż+B�늫�p�
��L-�GaZ��T0$���? .�w||Շة�ͣ�S��Lk:$�|���)SL| u+'�? ��:��ӏ��>v��M���ےa���Q��0nY�9�lBky'�G�Bg
4����i�2{�s���3
�����Uw���ȅ�,"ȕvE��`�(I��h�-��\�_�X0i���ܲ�9)�<�]R����������E�n��7O#��|��1�2υ-�Q\�����C�7�ڎ�"��D�	iB��]lO�۱���ǂA�9i�i��=9VY32tO\$=�����'�R1���z�(��T6�V~���O�����8 ���T�+�v����7ʣ�) ��r��/o�3� ����c�՜qzCI���b��m��7�n�-w�F�}F:R��^BH�zc�ꥅ��q�Cr��|R	_��1�4j�^���iK `�����]0��<#�'��E>�A��'��&ȗ_�ۥ����	Ԟ�"��QD��t;Xd&o�4��v�V�	���&q��6k�H��o���6Õ�n�D5m�)�j�1ץ]�~�ך��d�81� �f5�^�*\�m�$��DY�Ό�?f4 vQ��E6Z��߉LGzbqL�te�b���SϹ�e��;n��o[�8K��`�T�T��k�+��zR�>���k1�{.�q�B��_贘�wW�<�87�{�72�٪^�X�&؉�70B^��,v0���Ikj�Jm�	#��60Ŧ%��W����k���1�������{��{��[�q�[#`J(�io�y�;=�s�M��H��=9�� '���@���$��LO�4"��O��)S�H۫�nҀ�������0�K�M��RI�w�I�<"ԏ:YO>�Rx�gє��/�L�rلe0��1�A�d8���G�h�[�!Pb�j>���C,��[�w�����oGf"A��i8����n�<�C�	+����8h���3thK���x�p�P�J��OV�;�6Ԑ������m-�ş��om�_��nÏD�@i
�l�_w]=ә���[��i���_�1�HLū��KV.�����>�À�ai<�c�>�vϩ�K��ń�,�אV��f�J������.~>=��+:�L:�Z+�Ѱ�e�*��xۓ1�����6	
W�!E�U'�
���b��qNI��]�e�A�68Y1#�=`Ijk�9N�~+���u�U�f�9�ڀt;�FXV��.�u���h ��Um
`W"/J�U�S}�Iʎ�	�;£&�q�?�$ ԧ���
���o��goon�$��=V� ����{�Ԗr����"J2���n���gy!� �" �Z�{� ���D~ZG���\���R
X~���N=��q]fB�s�p��HH�j�S���=���d����SK��`����B�q#�}�VZ������Y̋���  ���`�7�%l̭�Q���c�i0�l^��i�4"�{;y.��N���jCX6�;�׾l��by��Z8|��е���i��r�o�&�󙨝�����[�=�Ph���b7���y�R��ǌ~\!c�����k���J�V<�!�aDp���";F�e/t�R���<%���#�s�
�ٸA��J��Rq����Cw��� �|��:f-%-�����v��L׫�8������ {ӅH�y�z.�&��D�}����I�ζ��Ho;B�����^�F1�xۭ��X�9wd	*~�W9r��1R�C�=08����,��s��Ln/�I\������bNpB~��*Hl� \�2w�B	zu���[^r�;��ad�F��Mך9V+bE���y杧%휹��e\��@y���"6��~e��H|����BY�73M�z�@��u�}�$䕲�=%��kxj�!��hd��ˣf!�9���j��[u)��)c�G�l!��Y�ŉ!�v�#zMG{�N�E+�� Pkk~��I���QoDk\�d��q�/��L�E����Οdg~r�ǳ�� /�r�B��eر���aB'[r�I�;��>���e��u-,-����?$�~�f�Y��^E�� L��fd�5��  )@6٘�����'��e�G�\�aJ\M����pv�"�]�󹓱0��9�<��zl$�f�ʟ�P�@��<�� ��{g��� �"R�߹������7�����o�B�w����0C9�+��݇��2[7X%����g���63`��ꇗ0N�Kv6�<\nԦ)��0
]�jS���Tyؒs��%���UU��*.�ݔi&�J�A�)��Y���why%�4?�͞�2\�fjb3���{@:�L�lo`G)o6�?%� x�W{�Bb��6�O���S|+�������Rk;��_��\���f���Z9��[/]�K�c���(M��S�R1§���P^8��������:^|yfZF	v-�2JK�����#�fc��!���Z9��J�S�4�����6��/r��s]�Lƒ��GC!�:K����_�&v4F���U�#+h<�`H�w!�o4�=(|�j-U����"���NH�6�C���4LQ�TܓE˃]����j?"��d�v˿�xc��e2�7~~�b��3˨œ�>p��v������w������N�Aht��,�d���;2O�^��޿�W!՝X�j��{})�B�p>���3���6��X�V�g*���k9~U�����h��4������n�^ƺ�=Mkh����ʱ	zb�U����d�w=[� �]4^�]�%PL��@�[Lio8g�_w�\`8ÀB}��G��:kvb��$�Y(De���E����Vk��?F�s��Yӊz�����Լ�^[����u�rwl�&�$]H��s[�c�����<2_9L[/u�7+JBJ$uԇ�u��,е��f e��I ���C�Θ��-�e��8�ɇ)�:c0�v��Fr�m1±J����a��>/�y�(PU̜oCQ�z/���_\c�xV#r�5o�v�j8-�5�t�BY.�o�I�����>:��jS6�#*��;��BG�3���!�؏�W9���������l��t�0�Nw2�s@Oυ�4�k�ԍ��y+@ �������d��bp	W:G$A�oK���L����C��E��.2\��>).��|:�MVU���g�|����t{,��8�pʾ�d���d}�̈��Ѝ��1�H}���B�?�6� "l|�z���璅v���.�$'�����8JNB�~56aK�[lkN_X?;�,��%!gx<i۝�'Ӑ?�7�n���WDt -�0��Z��d�! H�����N�PM'�JR@��lE�\ s�8'#�X��Vq1�q�Y�Ѐ�5x�rSE�����y$"
��}�I2�,�+V���4I�P���e��uL�����07�[%Ĉ���xN�CY�?�y�v��sl�R��ʬ�pG���'x4qg��5�m �6��lK_�^R���p�^2�u�
���:����%o;�o�G�\��k^�<Cx���u��`������z!�m�;4ô�j���v]	c�k�dP�i@�����D���QQ�c���%v�!(}�\.�[.B��SI�	=4��Ht��gH��^`��~e��ޝ���p;�(W(���{��M>� �Ӓ�f��@I��CY��L$,LR`�yw�����p���@ypY�a)���:'�tȅ}�aT�?=��0��̉�� ,�M�[ �����bZ����y�/i���T�Qݔ����f�j}�$�����\��	��&��e�7.�O����� ��DQ��t�tUbB �6�	�����6OދەS]CS�[~�ր��Z��5i���@���
%�AK@�P���u'��[�1*ģ
�t���Z��\��2��6�8R���E�~�c�/T�:Dss�~��Rĕ�+��
Բ�����	g���L;._6�#F86�-n�s�����cy'>7������Y�RN���I�0��&}S��oK'ΙV�}+|�bK�+�$�a���Å�W7��R�1_�u�cƳ:�(�ԋ�E��N 
 ������9d����4��Y'��/�ϿG�,=`����T�ҫ�]����"IE�]_P������+��,o�M+��J��g�9��;��?�$<���n�2�Dَ�@���~��aU�B��Qe����{���n 7�բ�r������9Iud`�rb��܅����VX�ao[RxJ��p�:J��*�*0v�����$W��
�?�h�K�68�^m&�V���P�ۢm��ά�#��N�n��jX"Qwc�����}��������ҹQ{Џ�.wb�Ԥ�$�$>��z�{��m�;E\wӓ�Z�N�t;J����F���ƀ�~VH\p��f]�f��sv��Y&�o�V�����JZL�C�z=oQ�MD�i,��ΠxrCx���^����^��n"�}o�n��4��e�u�9F�� ���ACQ�B M�Z�t�}l5;��\;�7<�Y+�K��I�:�а�-3D1v=�N�Y��?+�������hN���Czs��I\:�X�m�}
���>�z�)Lz�,6/(
��*��|�H�~6�,Q�t��D7�QTK �;o���>	��>�Xr���� �W@���^3A(0J=��� n��o�O3���-� ^��od",!z����=�<I&�B���?�j��n��\ƈe����S*��52N�3Tk`���
�*A�q�$����(���#	t5�.�U�Ċ����[��%��ѿ����T��"�0h���#G��H�ɍH���G�Mq�|2�L �. �o��3��#-TJ���V��K����\�׋��Ewݪ��N+�UIoʇ�~h�����JQ�WZ9�@	.>��WʐFB�!i,�g�铹@?:�4�5ٗf�aΩ7mw�h l�Z��.r+Cn��	�[޶��!�o��+7%@*�J�E���e8�gu-����ht�5��|�e�o��Ѫ�2��|F� ����Y�K����r�g�����rk�Ƨ�\�?���1dӯ��L�|K{@ ��a�0��虡�*}Kv��#�R6{�?l'qGa�k�"ذ����ؒ��S9BG�9�n�~�g��[w|�n��!�@��9w%8`S�g�Z�Ӏav���f|\q��G�����#¨�E�s��/o0s}a�l��
簨dK�{"3�&\����ca�x���G�7�++���Ek#e��\�G�n�u�ڼ�#��P�����7�L_��@|���D�� 3U�$=	U�҅��]�8R-L��O�g�AH��@�FT��>S�`to�U�C��
 �V�z���C]KkN���	�)�>��-4#a���"�wR�my�W�nIW�,f�K��8�������S�m�"�P�0[{+X*�U��a�G� ��?�$��N�?�%�$E��C�K-�p�X�����x����妷�C�W"6��� �]m
������/� �ML�絈���J�I���C�G!�<<��hŨ2i�.]��#�+����m����l�v�W��DJvę�Y��q��#5u��O�=���/��d��
M�ww[���^1}}�6H�ߕ��G��Ӣ�v�hu�r�ku�8�!����zL�M!qOuŞ�&YGAf7��a�	�P�h�[	@��y,�H �\�=5�Ż8u0}���)^�Q��|�k(R�r���Nc]�dP�i�M�wъݎ��)z:�.@qT�qH"e���i���~�c�_ے���>��
p��Iҵo�h��B1k����ПHYN�����i�R_M-BȆ^�̢)HRa�OZ˴ѳD2��2[;����7�g=�z�:�?��-3�lʸ>����F.�������	���V3JW�~�i�u�B��o�X�6���У�Ou��b/�@mϑ.��|�熉�Њ@*�����:O��d��B5��L���[�h0%���D:�ܛ�[�SDh������'cPx�����c_;=	\�5����C&9�!�^�����nOr��®�T:�S�ɴ�S3d����<5��� *���u򝤸�D��Bn��J���&�u�}X�/Mz�q�8d1>�$�`E��,�x@/�cq�(
l#VA�ʆ$���0��Y����!+�{G�r�ߵ6Bɖep��6:!ҁ�oIH㚿{�1$V�dx�s䯪$�|����0���uS�ƣe/�ӫ�5:�t݆� ���ZnVͷG�Nޑ_�p�d������Z���
ϓv?^���2�q�P��1����u�u�	�Z�	K�*��K�\H�:i��,4���<F��%9���ٌtH�d+V�>R�Ί�!��PV�����T��\��LB�5x�}	���)��OjČq!ԑ�z��Pӱ�X!Fk`ć^�R$:��r�uT�$aV�X؎�b�ڛ�1��/�C]a�6���L����@6խ5x� i�g�=J酔7#�0�E�������}���8I'�$=�<��雸m껯TD�V �d��n���{^e^���Ќ(�J��
I�}��7ʢb	&U�T�N�&����n���8�p\�	��)]�t�"�i�ޱ�G����X +�b?pD|�f*�y�V��k�,���t�[�>��Ba�J�í�M�G��8
k^l�^�t���;w_���ꮦ�?e-U[����$��WG����#|m�$M:��g���g���Ǒ�6��3(z��;�΍^�K���&�n�$���U�a���/�N�ˮȭ�����A�7x-�~��$���~Kt�)�0��8Ju�d$f*@Z��۩����Jn�!nr"�&Q�6�|��Y :�J�v�p�7t�qEl����z���Am:���d�d����\���t�6�P��$�Ҵ�-��- &c�Gn@�5l�0�G�~A>U���m��6����WH�O`D�.���'�W�Wu�(��<��u������]�*�.������@w��Yp���1&���[��;�𙳸T���BW=$�_7���n�a�s���h���W��A������$��i*e+������|I��kK)g��9�9�鵟�}#�FC����2�:��X 2��^�3Ӝ����y�r;�i�}�î���4 ���
�O�B]��&)~ef��<�8���e=jk�c�*5\T��׬�x�c���@�ډ�$��y"d��0́�m��0: 9x�n��,��ō�9|@"R��MU(C�w�p2(p�t�(��y��Շ�2@D����sO&6B8�E�Y������96ے�m���������j�P��'�=P`���1i���׫c~��|�RF���'��o(�_��X=PF?��c�yޢ�AV��X�+��J���O¾	��s�R\H�����H<�f�F\�Z�Z�c	@���M.O]�CR̈́W����s� #KL^�c��U���Xl�� �{���$ך�!���Bwb[��<��*�P:.��<l:l��&��
wًʹ�����\ug/��P�cd�4{d�/x%�~o��е��"��x�Q�����e�@q�i����ō�j��N����M���N�B�5�9b��Į��J��3{O���f�ͱP�j�(��f�*����?'�L*w�H�$�X<��?X�c0ELpt'�fcHR8^4;�q�C9�Gx��y�n(ŌV�-,Qo�שіS G�m�1��Ǿ�m��$�������ҁBΓ��dU�(�qR9z$�7�bH��G�5�'|��#�J�b�?Z흱a)J�鶰n�x�[�ғ Y���w��_�F�%Xa���$q�i�ɑ��y_��L`
ĉ�r.x�(�z����R �%�3���e�3W7���Iu8������A�l�5�C��DO��v֤]&�#}����K]:^�~M��Q��	
���)(�xʃ�<���.V�ι�-^B�f��N�M�;���n4� ��y���-˕D��M�r�mAb�>�.nl2�T����t���ޭD���N��N���k�p:��41�� ZM7�KkK9FM�;����ŖI���((�ӂ��f9]�sքd�}&v�6�D��ct,�3(�p�J�)T�a�|�u�g�.�C���]I�wn�� �9��謰ou�'oQ{�}��N��/�Z�*|��`�< Jr�T�;�rE+(�3�ce�'�\b/�m=(�^8������4�̈́���L�AK�/*d�P�&�ң���x�]�&��t"sJ�ELY��xW�t����\�žϩ���f�S�&����5�u�_�VQNO�%�Oj�����g�*�#/G�*x=�f]���&�bb�x�4�̋��.�{wI�����;�O;�&&�}�t�:����b�i�_/��@7[i(�l�/�z��3��7��edgh[m�!�YMGs�,<�ϲu�Gu�<�����ʅ�^��n.���r����WͶ��{��wj3�+��9)��s�h�!/^�'�|K����/qǰ�;�����=��z!UEB�qR�I��D�ܟh2Ra'�(j?�?������~�i0`��F�+ӉC������AA��y�C+:9��U��V���P�57���W��
���xEVU��]�&�Mژ���܊��DT92�y�{M����`m�A�uQ&\�1����k��
�	��q{�B�b��x���e/6��9!׳6��4AX�/2l+\'}<h1��.Ti�_�7�;<�� �^DL�*K:Xej���¯&�X/��wqB��^mk�S-��tF�I�-�4������.<���'��ʫ0���ka&�^{~���@��>�ͱ�x�p��c�4`�b���f�,g�?H��Xy7�0�.{q�@(�{��4��*-��^�P�(��^3=J�u`�ʜV��ND�6i 5��$�PL$ [��-�%m�|��N����?#/�?�	�B�{[ux�	c�CSՑ5Fb<e�`�8���ޙT�!2��ϛ��J-�~�(��x��~��P�&�'��x�����4�چK��'��_t � �a-Q���1�2b��j�[�z7�cيWv����R��_�*�-�>�2�؄_W
�R,�S=�'ˠtV��~S��eC��~7��M�vfA�r��Ϸ+�n��i��Mj��p�a�k���������G6)^zV��|��<ņ�B�f �=�b4N�?z��?�U�:&�A�[�
��F8t'A�F�_�ׇd�/�w%zV�PQc��aӁ2/���e���{[�D���*��l^�qK"��5م���j���b��j�5p
�p�	oj�
-�|s���7���n����Y��Z��{��0�c�Nf�$�੟�g5%�v���b���9�Х�6zl!�gD��U�P�1 �6.q����~��e������4��W�o�o!cHI��5S��E��o;����o�r�l��c����)�wU[P�7�<�7�Y�,�p��Z!�a���a�F�_����1ai�f��~◷�e.���!����J�/��v�Qt@�?i��훽�E�l!�Y3���p�;S�p:?�P":Ȼi����ʨ
w���jM3��Q>�%ͦ����<B�C<���n	i��&6�<f��>���G���e=Ƿv�����L���g6[Mz���<�!�������D��~�i����_�yi��(T�L��i�y|�����������q�(|Ya3K�va�}"L݃����?��Gߎ�N����E�%�l��g5��0�cY�^�X�nz �ZȾ���,�x�<�w����B��V�� 4�9g�I����b��pc��:����?Z�f��7��L=�T*>�#"�F9��`Օ%]K:��:	��}�2w�]wQ2�����}���0M܏��e^���b[˒5�0a��R@�l��!����VuP	w��N�i��C����׼t_?׽%|N]�-��L��TIk�9EF�X�ܓq�P�^�!�RPh����.��'�C NB�:����WG��,?#�����P��m�aj9T�sd�g^i2×�B1JQ׀�j���6�u���QTR��VA���$>U[���x�}w��_�TEj��	�����Mi䀲x�d�?��r�b��迡�_�(T���W k��H;n����ۢ�Ի��� ��J�Eڏ��{d�)L�9��7O*(ݩ�6�@mS��'��յ �o.�F��| �>P�)�4\�E��+�Um/���i�и���3�\�.m�L�x�����!����r�uJO25�p�Ӹ�p���
�ވT�2$*�t��(��#vʞ�(�*)	u"���o�i�>�F0Xӝ�^WrGl�������W���#w������zC�-Q�_5[@�v�V�`��IV_�qG���نC"�l��0b|��Z#p�$|����̓�3u�u����˨2����Fٿݭ�v�Ӡl��|����~`Dk�,��g3�B][yb;R]9n+7:ދ�K�n$��mO�X��o,�N\��5D ���d���wV����z�����8v� �L`�G�A��N��"�)��3+��0M������yÃ_����	��<KM�1�I��A�	��m�c,w���$	ч4��18p#�SW�g���0�ii��>�*8���7m�}�Vч~�o\���m@c���WC����n�}��>mL�Z����¦B�����D��)Ԫ�c�d��TQ���S���v��⢑b/g+p.}�|�6eoAbc�R�	�M���D¦nN�~����?�`�QA��ї���f�Q��kK����Ic�j�T������
�d��Ȟ����ugAs+���9#��:v�. �,U.�$l���r�� ��q��q'�s��n!g�&(Q��~����!��ޡ4�tW_��iq��Q��P��3u�)i�]P<��8���rc�I���c`����	� $&3Kv��:Q�9�o'���@X9���;F'���N}a�$�j��7�3]�om��p��!Qf�dnmzY�a�<~K�ł��,�U>��N�'Iب>�(^M��	)l,7����T��\���c`����� ����x�ٶ�I����=�?�Z�9;��w7��-a�5��}��B�_�Y���w���Ͻ
�����ss�BT�`e�i�
�^er�(U�O-��9�����=�ޱͯ�/$�Fh'w�gS��@��B��R)�~0�� ���a��%���[	
�jd�ϓi���G>nq�Y��k��CU�����[�����N'���묉s�{�R7�3-�u�O�gk����'��S
n6 �f/����?�ϊǔ`H�8�0R�y=�,��s��(e�O�*�m-���eҒ !��GU�fU��~E��d�p7�7&/��ۅو�RD�!xs�t����iܳ�B�����e�P\�z�?e|�X�j��1��.u-u_�X4�c�xmz�Љ�u�<�$YD�칗 ��8�.ml-�U��[�~V�}�`wL$�Ȏ�.Y\m4�����`�5���k���HwU#L��$��T��%@˚���L�l��&��\%X� �:qU���|�HIF�����`����5'��8ńtƱ49�g�����Zױ�<"i��SŶ+�UזH��f�tT����[߼izX��߯%�ݘ��r�9ͬѠ.7�.6��3�J6�Q�g�EL��ZY�LG����+�DNG�r�ے�Z|�H~��:jt���t��Ƙo`A�0L<���>�(�p�Xu�˜�:zH�Xg&~��p���\%W5c���!~�I��ݵ�f��/,~Y��W��F�4�)�2r���@�-�g�"H}R�އ�s�Zt�^��r������徙N?�[�T�U��u�$�D�����dL��N�W4D�6���9��M�5/��'�����w�+=��O�ݽ��Q���U�y�ߊYA����������V�F��Uv'�a�_����aH��B]�p��$���0��O���rh�̅]���ǫb�� }1� �(��FT�:��+���a}6FS�ɻ���|ٔ��AQ~�;�wK��|��3����}�D� lT%�R��EW�ï0�[�-e� ms/�ʖZ�2�Rd��}�%��L�[ͫ�%S�;u}᝟�����I]ik$���H� Dvp�.�cr�.1
$6I��n��Wy�����KMp��s�|�V@��I8j�Ɠ�����䛖���$#�8���z[�VCB5%�]_c$ .٣�Vaכt�9�(B���V9^�X���Y�ۮh/
�R��K�H�l��q(ſv��>��/��ɹ��mmH����I^���#�ҼӨ�'\�k��0�n�BՁ�~�����\.BX�� lX#˔_�O}��H��~�PQ~Y.���J_�ឯz�UfS�����c�yH����E�:N&�&h���>�oDD����t8��)�r}�^�T�/5��Ǥȕ?:/[s��#J��+�DRH����x�量�N_̷��CC��7�(�V\u�!S�s_ ��K�%���84ˠ�f��T�FǑ����15}6 �	�zNmx��aͣ�_�r}�!�	B\.�:p� 
y X���u���7��v�$��^�`���e�����T�I[�-l�� H>�ðW����a�r ���c�(@*~X$ϝ�|5XN��맂��dД�e4���bL[3�-�
Z�p��1����S}�&)���f�e�#>�]�t,>��&��}���q<�Ma𥃾�g.�"�����mi�|7 |�o'�j�5}��'TR�<����BV�N���<�>K�p<�lf8�B�k1'�3;U�_܍o���M&��J�C[���&�f�L��̎�v9[ڷ�*iJ������80XM#
{Q�@���%�c������ܪ�{@�ͤ���X���{鯤O>�h�8�}c��=Q���˨���y$Q"���6
cZ? x`�����u��#̡=�[!i7�2��A��"���1�#_l�~��;��yH�g���",�U�j��7���t�J�GI�ƀ����K��^��Y{`c��C�-76��?��NȥfM�(���NmQ\�G#"=o�z'hOv�ӵ��7U^O��M����1"+�a��W��-D��r߸�m�$�U��^�v(�����7;]'J`�3�/i���/���׋��K{5��w��T��)pF�p�_���Ze���ŝ�B�pM�P�<���Gꦌ��-��LC���%Tmφu@�+L�V��$'��NA�D&��2�I����0��!��	��uR�(J_�a�%��ёS�@���mB�)� ��&3�.��7H���LV'�G��,�K
���wז���f��%��Y����a�m���c����v_g��<�����,R�&[|�qD<�M�è��KR���4�/L�7h8L�{���P�m�~�z�{�w`F�q�۔�:��g{�#j̛��W� �M����Y�7��f�O; ki�{f>���C��	�W�&��zYi�\�2��}m�t�'.�k�"L��*�5H"xSW��w*�ܗ�.&Ó���8�v��B؋�r���d0�<sOG �!���(6h�;���7�O�G�p˷���<�����H?�#`��sk'h�;�s��$�1Vذ���q��<��@Ds	G>q����A�L΀;���cs�¡p ;ʹ�@����R�v�����=���u	��x(h���M��>rp�3���~�5I�g��.����K�4`� O0hA-)t	d7�>JHPI�ϫ�3���Pb�
k�%O�˿v�	��ThX�@�h����p��)�Qsy��0�hD�m�#�;i��C�VH��X��5Y�hDҎ�C*��4�6��,��Z�a������Y�#lN�_E0���*�c�Q�ΓP��>pq)U��=�E_�y�BQ�xo����"L�D�x!f��dϞ�!5-X3^�{��T*v�Y����=��6����r|�4��|���^/ּW2F���[ټ�����S7G���s����R��B��^�R�i���dڲ�%g]�I��*n��H'�'g#���9V�������piҗ�.No�z��1��M��w�A���(yU���Ge��� ��/���fO,u��5�C�zq�CHAg�'�/���n�:`��U�yn��=5{�0ɽ:��h��U��<��Q��VÝ��pG�y"�'��{n���J��+2�[H�<g ���'�snk����I��cQ�˹SA�t*�gY�g�}�W9�O�6Ly�df��*D :a/Z0�c1߄m~��g����d1�p¶c�=��VK/\��\��{�;����9_\���$�-�Zh��	(�uF$k&�
v��A��c�����0M�G�[]�q^�BS�m�<>٢K-nE�L������q��<�0�~<�\�^8����.{p���M�~$��9�P�C扶�^t7�Ϗ���9.�����󑡩����ao�S����/Z�މ�@�MT��]�������M�B���C	��?=@F¾��~�� �J-ob����CɌ���W$�a���肩:�/�����G=_)(���n��T�j��j_�����BmѵZ������q�����Jˊz��Xͭ�.y�:�j.,��Y��q	�W� �[w\�c�5`���3����Lxd0_��Hg��}\I��z���dņ�� 7��hrɥ�7��>���7/�Ȅ[�kEv��w���e��7��CG>��*�YWF-0*�ّ�w#2���H۔%�ǖ=�ٲ۬�Czh�xNBڙ!^�������=�4W��\C;����jM��Ea���Y'��:\�O��ϲJ��$7�p�ը@�s��1����w7&�ME�9U�/E(�l�7����3z��#��,~�J��Ɏ��< <�:g��Gإ%�#<o����JQ�$�J��,i�{���kڔ�?�5;X�{m
��YU2����|����%-����W�[������0�p���¥��'�J�lM�9G��e�?�x��^�,X�v�8�[?��a[d�bm�2�K�5�Ҟ���V(�AI�10R�D�q�~����L�}Z�A�7�Qk<��@�4h�|r�����A��5r����C�$xZ$�%2��~ ?#[f8i����tW��wx�ݶ�"a���hٹ6���r�U�O�1���9uobJ�Ӟ9͇g)���������#���Zp������l��W��Hhy��bwOs�G6��%�X��ZW���/!��u�?�d�m�>6����!�I��y,r��m�"��L`Q�O�~ Άܯ�*�7��?K�I��m�|@n�d{ ��A�N-Ӎ}{M����Ï�>�~�Ko�O	3���:��!�R�q��5�y�4����ʇZTA�*�v��� �bk�̚��P�ʧv�7.N��0|�@�:������=�t������Q6��E!i��i��w���U��^�'0� ��k��;p�5M��B6̙J�q
kb;������x�:Kb���z0 �o�kjJV��m��v6rБO��Q>�vr<���,C�/� ����뵛-�<���<p#sL!�dX_˦�����mT���k_����U⻄��ٲ�l���W�-�5��#g�e�����g0J���&�8h���
"�ve~�!���0�0����ODΈڕ�oGR�����ō�0�б���򝞇2���oUV!��7](T
�7"<����������x�<ց��I���F��6�a1�{h���=���Ͽ��"^E�<���G,Z���#|m �Az�I)Z^F.�؞���L��{�P��o��MO��2#3��4y��H�K�������JQz��[�F6��8��OXԡ_a6�ή�bC�$j�A���c(��;$G�IK_Y�l���\H�9y��H�ym�Of��FcF�v�#hĶ��� �Z�e_���rAO/�x4.������I1��j�T�Bî�Ma���f��"#��0
�G��8\�b)H9��p����-��ή�/@2H���A�k��z��N�P��7v��I.
W����|�"+���|Hl�y^����I$(�]�Ӕ�~e�ͫ�����Sh���Pv��6aU�Ice��eD�sb�|ΖL+��̹�/x� \�c�<般�>�X��.r�z=��oh8�a���^�$��������5�g~���q�@���`���9X�m��}B/���u�P�'�J�`�ٮ=jrS��!��<=1m��v:lM���YF��% z���C��>�skIsZ���`��l�䯒�?��nZ�+�I�͖� �s�7&�0nX�*����M����<���d�v]��hQ}+�8�qA`[�S;f̽�����w��s���ʩ����_�l���)���	��x%�����VV>Ҕ�%��[Jk~��kz��Z���k��z��4�b"i0��(��.�%6�]�[D�h����#=�����������W̰���k3���{��H$@�2+��F�N�,�`3����hg��x��"�}���&����gއ&MK%"\h��/zI�w-Cyj+�� ��M�#�c��߿�F�*�xk�\��R����P^�p��?[�P|ȿ4�l`�d0��w��(��ɡn�@�w��W:lma�L�X���f���x�%囮PUQ���5l����( �j6��9�Qm�+ߨ��QL#K��7���}����z��K�j1�iIc�4|N��M���ys��Z�����$ȧ�[K)ɳ��{����<rţ��XE�>��wl`�/9xֳ:(�KL�1��C?��~�S�\�������J�����6�w#�S�!ՃhsO����b�0v�I�2��7��6��*��P곾�P�xw1R�j�|�Dp��&o�}�I�W����nA �W�z�i��"����#E��5��u�m��>s��X�;zR��6�M61��T�!W�<~A�ms����E΂Bu��!io��s�����Nh�p����J��E��������eyu<�H��/ť9\M���}�Ԁ�ǭ��ե�^	z��Ob�����#.�e��2 :9T���)@9�� ��R�1��-�ä�G�KJ�(JLn���h���,�̱*e"W	i:��x���7s�
F+>^�L}�#�y a;�P�U:��jq\�ad���!�aO�3���m��I+����M�*��݌Q���eԐ��b�Ft	<XV��	,���_V~�@�|g����o]��w4&u�Ac��O����p^p�R�����h?�h�"U�H��H,��l�U���7HxOݔ��G���!�kJ3��b�+�b/���6L?n6��YG����q�f�$�V�a�sG8���
9�]`~����^;�<������*��W��7�K��61	����~$���F
�*���y!��6X�ݎ��( U+�Jt�5	���9/z&ؤc��u͢T�Vۆ�*��Bh��h��*i2��1��ٖ��
 �.��$ō�:��o��9G :�7"���B��=� ��_s%Z�쌅ܪ�$b��������I*-0{l2q�������Gh�Ns�=��2{rV>�� hm��%Tؓ��*#E��D�r2��O�R����L!>�[�K�Tk��|���k�I4�q}A��q�63�aWXJI�s���t��NJ����I�n�j�� *YK�����]N�<	з�|r.w��$&$L����zI;��i�W#�IP�����!��9��ݯ�f!|���h3�޴oU�Tq��4du#��`Blؤ�a�؎��&]�	36M���������a�Gk`7$�o&F]� �}�ƣ�O~���$L}���2�f��j�AJ%1%GhU(�0tv����*tBO�H&<�d�B8G�XVN��)��0��7���~��=�g��?Q����'C{$Eټkj�	�c�����V�f�F��}pcÑ.�)W�n��I��;�=5���ar�g)+�^����Nd�%��'��Y�����6v���~L� ���ׄ�>4e��"X�ҵv�?���jMq^�F���H��~��u7UB�� N�x��4г�ĜgƆ�:�?J�_��]�[/5KS��L=����/��$)���O,�{t�f.�5]�Z�h�|��,)�^�HY��R��6�C8Q3qfR��KR�<�_g��l�"�4��1��T�.Ã7�K�̕�L����煝v���d�Ыr��#�=�c���M�[�E/�3`���9��C2<��O�0���s[� ��u�6���9�Jܰ�q_����"�j��gB�;^�cmuc%[.���s��%����>�\��$X��4�^����W�7f0���F*�NR9���� Y�$f��'z�
?�SH+i-�Ά�j|����xz��O�а����$��xv���Yo����s ��?�e�TN<��N~~x�}�c9G+�6A����tТ0�6�ϛʼ�W����9%P�M�����Q��j;y\��ǧ��b�+�
���~{��ɖ�.��P�1�L��P���m����0�H�-J�!��ux*�kW�D2���WR����
�������:w�F;>T������7��&��R���&VK[���|��X�;�k�{VC���q�W�G������]�a� Щ���qНbHGeR`&[���ԩ�a� ?���4�K���9�W}�2e��ǧ�~�7����2d�+�r5��VԐG���)р�A�ye���M��l�h��5�e^r?B��o��"�Ƌ�m����"�{��a#�x|�����Y��?���T,����ݩ��x�*��3?CY�j�+yY��Qɶ{�'�3C����v�z��pw.���
֝W{=�z�����E���ߙH���7��,y�2��j��7K�TPB[��r��2�;�C"L��[6��	��=���:/����5��q����{�0���)���R�'�ܯ�8��P5z��< �����'�j�8�B�&��� p#(����t~�
��wvV#����`��'�U䒓�D����<���xݭ�%���z��)���U��݉RHy���hz3�}�`"Y�隝1�K�w4<ȭr>GEy'��Y)w[�,�XaJЌ��fu�ER_�ｇ������ԃ~�̶��t'VY@�FC8����d�ֲ"e=�w�# �h.������
��"�(,'��D�1�d?���ޚE�`���Ls��W!��?��H�|��>��'��������9���T�G��1ss���&j�>��M � ٖf֊�DOw.�
�B���Z=�x:�GىV��V��l�*�㼇i<\�m�1N�e�/ܜK��m����#�Px�"�#$��\�9�´g<O��Ϊ��4,�f�d(�����v᷊�V0��h>6�aB
y��k�=�z���2_�&��)��kK��j"
�[���!�WWSlnfۘ��SyUT�k�~�r�:��	Ƒ�@;!�S-��|��Sy�)x�Ni�C'1��ԙ�k�;�����L)������g�d�v �h�|����Ñ�4�2e�s ����2` lu&�B��/e�dT��Fy��'��^��zH�n����J�?�؝`�cM��� ��"BD� v�:`�W�9��m�� i����w����*�{'EW@�� ��,�Un?>
'�,)5Qc�vJdn>9D�;[�P�@�U᧜f��xe�;��� >6U)�Y��(�+)f}�1��]E� Et���?׺е�sR5U��5��ߴg��b�<q͞��G̚K;4��~���!�4ê�����n!�}-U���'��Ĵ;���ԉ@W(�)W>�����k��_���W�t'a��Q=�OQ�# �?\
.m`0b�c�>~�G��/��k�{��CY���Kt�	g8�����:�����ڀ����<�� �b��R��'.%���b�Ȭ8��4w�����b���s��X�u 3v?�|����q�$��ث2�E�ɶd3�4��\_WE�X0}�+ƥ}`M#�Vc�C#�Ŗr�������@���ތ`}̉+��^��U��m}XI?<U�lYE@-�H��zO�_��-�F��^��cp�bc
,��tk^|��c��+� C	�x�'��"v����n���a3^D���S?��1,3��]E
S�8Q���2�	���m��5=������,s���h��ly>y�@`ϯR����=�.t��P�!D�h<RWZ20m�]X6�w+x�GQ���/]�Ԍ�>�f�
�)T�I<�X�2��q�8e}D�[���\њ��rN3�'޵b�C���q̋ݜ,S1�Z��_u�'#s+�8�(�x�u=+���%��Sb�c`**_d!��?�
~��:�0%ʜ��1q��;0ab�dچj�{���r��*_�n�g�Tר��2=�-k�J���gI~0�cT����Η���=$�L��H��Ē���zH	,�MU,_�)�mϨ��X8��\܈��1f��&i^I�6Z��̭ʾ
�±��{N1H��J:�3��l!i7O�^ x�7�l��;U�."5�m(�U��K�A}/�*���u��
�&�$�ͩ�\�C�#�+ԇ�w���c=^v�V� flxR��ƀ��e�
6�o��#�/�-��4�=i�}�B%[諻����[}]&���&�"�p�2@!��h�ͧ��֎Uސ�[�����="�[��dx;DٖT0|��Dq�<)���B�&�$�x���%��a�	fπb���C��{�������]\�!s�J�a�\R&idn�.]��ԭ'X2��$�I�ѹs�OA�O��V�qv�@a�P��f��ޟ�	xB"6��4eǸ�ka������`�G]�L��.�w��[���Y�-.B@$<��\���.�x5�i�	�T�Wqv_�Q~Y��09���5p���7�8�ʸ�!�<�&p�H�)�414��d?Z�τ}�DNQr�1dK���G����+�գ|^�ɹ�ѻ��y�?�+a�b����-�mRª���9a����?�j�$�����w4A��gS��=i��e�����%��� �(j|	^����'ԻS�h����VJ]'!�]g&�'94�큙���\��A8!��R�|r�h-)����Y�� �Qk��B���r����yU�D�s�� ����Y<D��G��E�c�ĖU�е��yr����4�Փm��2�qV<c���n��㌀
·���@5-eT$nYމ�c��Ӗ��f^��]��,�T�*A��v@���(�)�Ǵ�OB��p0��YU��⌅� ,/#<UʅB���c��G��X_�eT'�MQk7B��	2tx����kR{"�����M�<��R��-r����^}���6w\��u��B����w��pG�G2�k$ �
j~�����*HX��693��=����~�g�4 �ѐ.2��6�2���={�ӈj?�E.}���mr'��@Y�"�>�Ā�'ش]�Q'sb��E�+�DK�Cͬ:?�}��鮉Lb�6��y�2l����
�h'�^�l]�f'�BO�Sx,J���m�!��$��Z)��V���4�aA�"��ٿѝ��H�R�9����MK�O�NU� ޸�!�a2��i�vȂ�BB98Ki$ã��b���E�y�������قO,�H8�,7��pM-_�>^*�����+H<4`�pt=b�3���K�q�����^glxY�i�G[d# O��%��|�^Ż@~�^/],�y˔n���7�U ��]hTO
��}�M��C|fx؜\�%�d>'��<�R��Q�syړ�ǂº�)�e&���v��O���#1�R�c<r8mHl�nzI��wAC��e&��7���tZLL[��s}&� ϓ�����wFY�R���p啂�=��:n��Zm��+|�~����a���������<NǛ0��V����:$"�*$	�]rJ\�/�H\��v�-�V9�fnm��ۥ���[~�i��ڶi��l]�۾��W$ ɝ�`�tlTB	/��V��f�:9:�(�芴=[���^�i��U-��{	��a���x������-����v��h;3�3\�5��"��l��΁-K���7�m�к8o�n���J �姕z\�	�j�����C	�[zMc���Ku�j��k���=7�ͥ9�������| l��e����R��p��"�\o�_]�Xr��3J�6�4��Ɣ��ͪ�]���~]����ڤ�����<�G$Q����pLh�<Q�����(��T�(�3 ���ؾ���}`H��JJl���k�r����iV�[^��G%��8�Mz�f۱3{�<��`����.�㌞>XhS���<"�*��y'h���&@$�L0��?�M�@�	����/So1k!"��Q��'C��q����d���f���E���`�|�O܍����<���z)[r��E����I�T̛������]���4�c��� '�m{o`"�F��o[��,1�AR��a��!�%��S�����	�L@�9�}w����zC����N���]m�|��E_�	qpl��iq��R����s�d�!,�Xw ��HrV9H&����i���)|��f
>�I0���^� (��;�/�k]R.w,���\�V�K��T�0����L��_��$��A��:u�^@��/au+\CG��c(Ҥ2���W!�U�$]�~�4hT�+9F�l��oV��3h��Q�%����~Y5�qW/	��Io� ?X`)�_�z� PN��گ���`�i�ۺ74h��G��@!Tމu�C�3M��\͏�"?���`�h,��ji�n��B�R��Yy��&�@0�ɱȡ��~��t�Kۜ��=���8 �x��'���a����+�8�t�}7�\���E���:���et�k �0���p:�1�H���-Y�u9�w��y/s8���c�1 �ڨpb)\�-�=��������1�t�i�� ��֞S��MI�b?��+�=�B��������?4�B���_8K귦'�_����(Y�I�@6��D�m��D�T��|8RO�A�ZĲ��������*�x�{i	uG 3Hݞ)%�|�yB��0��a���y����=�q�+ә�D�3b�J��,�Y�Bzf\!!��;�� ���m 'p�f�w�.zQ0=�@�e��T���L��E�)����tJ,�G�2��2�������3��.��81�NF�7=�f�7��Y�Rm)�մ8���L�i��~}�u�ee����/&U�kt�H����H� .J�#TB&���7��O��ڕ��U����1ʕ�V��(Ӭ��G&�@���g]?�q����xhq�l E�ʱԔ�b8��ɟ�R=���.cM@w& �-�/Edq %`/82g
7̖p�oJ�0�oN
_5��TI�߮�)]�)�ۂ���o�
��>4?"��#y��H�H#�r7!��(Jﳨ!,���O�/��?;���`�{��� >�_�B๱��� ~'�U�#��q�Id��"Fj6~��5��ǭ�� +:���螶:e9��z3q-�&�%+BǔL(/ʿ��]���� �q�2g�~f=^�	�n���P�R0;���`��h��v��&Q?gEBR���k���8�B�l�c���$�H�H�����ii/����2�iG�~g>��1Q�cZu"5ţ�zt_a^'���r��9��2�1\ĭ�x��.�;W�D��z#���W%R�c�c�����V��_s/2b�	�Ri*�O���<�����y8�뛂S%���ú��h��du>���+pPGQ��/�.Bd/a�unK��D״�X[��רiB�|�WD�맣��cU��n�ZEmW�b�o'uY�G�� ��!�|��䇈Fd��i�+t�5�T�aC��Y�|�T>V:[��
{y��y�8�f���EeL�XVc%���;P{�t&B����p=���6��	"]"G��\0�cyW%x�9�{.����/2�۳�
�ή�����{C��ƞ8{#��f�e�X�����j�j��jv�����u+�U1�
�`ކ[z�\�3G} E`Ĵ��� 8����r�j
��%�lz��
e��)a�k9�s�92֬�7��b��@t�;K���XY+(!z�M���h;�����/
#!㙥S������Okܠ�A���z��P�4��!%5?�/ϖ�ɉPS1��CԊ!��x�R�۝��'n�$+8�%|}��)�+�\���\eno2L�E��w&�Hwj�*�/Pl9:M�W��66�]�ܔx���gE�J8 �W	tH��k�D��bH)�/�0�>g��!��,Bط�	=*h��q3���Dh�f~SU����)+ '����y���>��Q]�m�^��S��v�X�8&V)��]��)ǭ#ݫ�D��J���c�Ѝ#x�����'Vӵ�Ok� $<���ca܃�<�̊�խ��z�Hk�T:GJL7���׊�硼�P;��K�41lr�Y�N[q���ּ}x����M]�Y�p�ÎV����.�}U_�vEH/� ��.�G/g�L2�����d���+;��M�/��t���k�)���ƫZ×Y�4"cg��� ���A޻\L�8�Ǚ���=�����AY5�u���`	{�ݫaP�[��$���]�p���6�!���ǉ�t]�y�P�	{5��AD�]<��Wݪ_>_�b���6[�g&L1tX�.Plspつ��ϯ�s�#8q�U�Ap������u��݅�y�ܕ�x�(�z��j��K�d��z8�IRB
#��{�����n,����N О��y���ţ�5�b��⛂��������w3UPw�tQ����L��,���{�t��� =@:|�����aŋ���U����H�t%���tR:A��֗�	���W�x� Yqj����ͧ���.a}g����r�l���-rн�k�~�[�����C(�H��m,����rW��S�z����&�Ʊ��Ã�� �)��XO��t��<���aG�O6Wz��P�4����ӈG��Ƚ���y��V�˄��x٨��S!��9/��x}��_mUR���E%�5��H�-�٤ĳ�ܤ�����Z�*!$="9�AԳ B�5�t,��l���I��z5��}����_�ۗ���h�?��f�S3�H%��M��B�)s� ��-R��%�e�۞�����Ž�������4�ޣ�m^�6<��r?`W���`�:}�,�^�\���j��J��#�Hr㱾��B<�xb�F���v	�"K���4��a;|��s�m��Ua�:ް��u4�9���_�G�Ȳ�E�r��/Xt�n�cQ�����S��>O�r@�"1/��������o��N�٦�rʾ3�/�/qrL0�����'�"����q�S��6dw�ׯB��ߍ�[�֖"$V�<9��@f��m�X����Č����{�$�ʓ�ԍ����H�P9YP���:��Uh�]�S@a ]K��:��Q@�a�w)s٧�]�#�Y�U�gQw*����@�i��B��];��o~��67wJ2͵�A�b��a���;8���`�ح����]�h�η��hdki&��غ��~0��蓦�����m�����\��X��`�/nhB���iR"�s��%�Kc~$�ւ-vԋ�
�����s���wop�a�w��h�9����ͳ�N怆��Z<ԩ�̵:NHS{sA�i`6��P��.��!vH��Ʃ�C�����emDm��F֑��ݫ�g�f���]��2h<�ڤ�(�L�@�H��KS�� �
	d�K�@�h����t@��*�A
@��7�&N� 	�j��뭁B��ߑ�l	�e����̥I�̀>)���.x7��ԫe2aJ&x$K��1�e�Ȏ�V�)��1\��,�xM���1�=��
s��<�-ՈS��篡K���_�US7hZ)Ͼ��?�:܀tn#r���q)3W����H��֫PYı�T�q�yi�,�)�A�ȵ�y8�3�8v��r��m��^����OP�z꡼zC�7c�zL��/��(�4+�']CGw|V�-�̓W��м��75r�-�K����Tj���=��Qw�X�I]��C�'���O��c���ù��ƈ��3�����l�5 }�V;U{����l����"�Y�J�� +^
�K�.�o����*ze�$�o,c��1��}V�h�n {��}�	H��r4��q�y������R�\߭0��n
�cTmy-f�����5L���u����]΢}�%2�XEŎ�em��}��"�D��*D���DYp@&x�����������״ #��o $��i1b�N��@����U�.r�D�k9��\G��>�6"���!b@��lu�Hi'9�t�����l�G��B��M��OCź���J�-�k��u>(�*b$�㣠�R�<WU�MV�]��p�;X�ȏ~�H��Z�D��a�Q�~~�X��H�������s�����Z�Igw;` #v���]�W�1��l���D/&)W�"�����TD�E�����*�����Љ9�������Z9�ܴՋ&��d8�O=iL�
���*� �����-��wg~�ǋл��+c��AM�fy���ɣ2�ج��j�F#`����q!/��UK�&����0����j�Z��T����H��P�H��A9rzӬ�0#�����T�)����
�$K�Z�0������6cf�M�WFhp1Y�K.�4r�Ԗ� ��B�������;�O\���:��*�CS��4�d,�Y�m}W�� EZ���ס�k��,]A��*w��� �mva��Of;�̍T����x��3rކF9-
�5�;'܍>[�~2���~%�B�I/������48�	V̍��W[l��6��B��$�2�d�r���8��x�h�zEYԽʽCz�����2�i1�@�����-��;����z�_0�VU�;��|j��,���D�z*P���n���g��dn��v���O�U���D��uM��m�z]�+�������"}�V�=�H�����w��N?	�}U.(j�>�� 4��� �/�H*ce��3��|����DsSq�Y����q�Kob��!�l�%xy�l�[XV��	�.�_^�gp���"Pfr4+8A�y�hvCȞˏ[���
>�VUݏn�­j���y��B.�<�������WР-�yF6�A��1k��X�<so��K�h�;�[�|v�O-�v����HJp��AV��U���>�js���n7�D,��I�O���t܅eZ��i�śG�_AMw�&��=���1a�D���*I��^ Z����p���m���~�M��zC�,c�6E����MBK|g�[O��B�$_���Q`���\�����l�U�� {�l�'/�N��A?� ��I��i%XN���e��jQ~w�Nwm�⋙f �J������\�P���n�g��[�-����[�3c1?��`�M���u��/�$g�/��Й��qT���i����L����dR�dO�,s�M�@L.FM!N۵�[6ݓ@ֽd���ű�l��&��`�� 81W*�ZWV��T>���̈��w�١f$�~�?�V�c#su��g�mB�ӳ*�����2:� ���
D�X�\��,���x	 �h2Z 
�~��8��� >�#t-���З�B�O:�&F� �Yok%l������V�z?cә'��LGє0ۙ���42؉0�{O�OPM�������3�CE	��� 1�u*d*�X��
�Q�2�a�۱�S^��&�5uȣ�]yh��h��1���?���BbK��Bѹ��p=/�@�����������$�i��Y��%)t��|�j�S1C��9�����C+G��Q�F�S6�	)�����t��gEà�;#�,�.��n�qx?1͝�η����t��6�Ekx3y�L'w�IZ1%��?����n܈?
�m��h��ູD��Y���iHi聁P6��)�V��� Pk#,uen���Ş�yS�Jbt�q�b��YZ�����bx��>w��B�&Hx��q��6IqO-��f=�wp0b�s��X]ۤ�[�H�̪��*�i{ȇ��i�+T�F�J�~�2�c�q�= f*����|�M��ؚ�p��!��>�&n�����k������W� N��j��V�N��-b0kۈ�����'�T+{��p��-��z����)?����&k���W��3ukxb~	_CE��M�m&,�����[ �w�qeܢ��sˤc��C��32�b��bø��z~p�~�6q٠*�uG�;��y;�	wa���`A��c���2��%��K
~{8s���^�^�s�-�����1�~8kuU3���C�r��݁� ,�~�G2�\-B9W��NV�C����;�Ahd�/��Q�>�i�챺�������Y,
�~���
t��_Rӌ޻1E,{�����_�܄�hPrᖞ�m�V�� �,� ;��PA�J{��s�XD���;�}��x �k���6�n[q��{��������.#��T��xbAZ�u�= K����(�_F��b,R��� �+Ghs��*�ё�1v�q�7�a8�3�%H���C=�-߮~��7���N*����������,dU \�`��!,A��E�_�b�bµ����%�Sգ�o��z���W�Y����:�ˀ�~�FHwB��	��J6��>��K'݉$�+t&�����
p_'��r�S7�{o@�G��(s|B�\�����"z��*�dx:&|`=����0�g�<�i4�P��×a��,ԾEL�)��>���oRM8Y�J���J�f���W5�!7_dӸ6�yɉ��F�X�b�N&�5�F4pe�R5&�j��US���Z�_���%�{7�1���İ�Ai<ڡ������1$��ܾ��HQNN�	�#eUo����{P� ��lIe����
",���c����*S��C��V�q��jc�
%��Ce^�4�f�E'�Fڙ��`nZlb5K���}�����/���x�u��O/�*�N��Q�+��%���R�����,���G���ak�?���MA
N�<�)T�6����t���6����=(�}��eS�]o�λ���`��[6�yխ'8��\��
(s��8!�E�Wvmۄ��$ĨV��?�=�D#�W��Vd�نQ��n�Wط^�O���x<�o�Ի-�o\�4��@�3�)�X������S��W'���ܰHW��z�/�O˨t���
�T)0���(��ۣ�6�Y@�&�F[�g�B�C�a�Wr�V�0�tL��������5��(�"���W�`�dU��1�5���\��!��|���� 7��G�@�a�j̄mK�?��,Ȫ��i��bs�5��T>�h22֧�|�@r��fN%�.����
GZ>\�v��	�,ƭ���t���E#|��-ɿ�������6`[l�-�.��� ܈�9��;x�>?^3|H��
)��]��O8���=�\�b|��&O��k����NV��'%a�v�pr�>� j5��a)l\�<i����+<P��
�Ƃ�-��6�b�+aŰqIe��ۏLt�sD�OTk�E�`1�$@��zx	8  �5���Qی�mv���U�3ߢrB�6�T����,T��ο��8S�$S|��6�@ƨ~��Q3��$Tr%�펿���Nثs�1W��m�E�1J���+h�ob�gﻵZA~�\"9q�[a�oTهJVs�\����F��^��Ś���L
ͷ������r�N�I���$��&|���!$fR&���=���#�d��O�
���E�jn]���b�V�4�A-+�������W?_ՠ��@'>���&7�9�[ϛ�6��~lL�x
?mW��$G�T*@0/1U�����yB�� �cG��D��K�K�|S�r���r@ι(�l�E�e``k~\�T�"(�����&�k�������{�Dם�u�᝵�֋�d�̽��?s�������Fr��B���j�(w0Y:	��Ъ?K!�v}�y�&��]ߕu�ߣ�R:LlDh��N�xL�~���4Y��ڊZ%Z��e�|W�K��\s�Oq^�������N}�4H�+E˫ޞ�w���: �T�g��d]B���Lƞ}�������Z�|��]�_ߌ}�H�xR?��BغL���I����%�z� �j\����Q��s��r
@��o���Km�0�����
���2B�W�������[>���9�?��K���b@2�����S_AH5�m�K�7�O��׽�`����q>y����,���U���$�a�sڧ컬�ކ�kq�tǅ�6G�� ����দ��k5*�g�H�d�ĉ[�ף��mEW�W���Շ�9OA�F�ҫ�@�i���b����*���8V�'�.3�[���)h���Z�,`����`{����n���A��u1�dT�/�=)5�K�Y�!K�D�hz�X��:`{�¨����c}�\�}h`��-���X����N����u���[�8�V�!��l��j��\>��J�̸�)(0M�o��/T��d5�Tg�{!��Mͤ�mI�b+�߈r��8]����H��|?��9���z���1�C��K���`�g���n��	t�=N'�:O�"}(�Q��d<6���?iƚ��r�.���~(�:�ϕ*�&�SVk�&j�����t8�`%�}�{ZY�h8=����Lp����⥺v�<r���w	�FF.�x�V��Lc��Z����q]��T��vi�pXnTٿ���A�ل�id�f�@s��d-}���u�<@Yࠆ4�B* p�6M~{���*�Sɖ�|'Y+x&y�վ�ʠу�+�'��[Zė��6��9%��)�W �E�|M�Á�]���(o#�\[��ה��X�������@�
'��P�|��:k=�W7�ƺ�����]'n@�e��*:�ِ"�����P��`���e�o���(��rn;�D���y\Zf�,�������t�V����x��I'�ZǓ`�1�"]�h_aո��E��&��/g#��d�-#D����80�o�a$5P�T�c� F���$���|�:k<Tp/�!��g�n��Sض�l�1�7Sk�Kޚ�p�[�a�b�#�n*6B9k��D���+7*^�[g1]���$J_ְN(�Si�Yvw~K�����XA0�e�!�>|M�pb���8p����Y���,3e�ȴ\���m"�v�<eN�y�B$��h��Z�8A���[�7�]@�5��v�|g@Ab_=�w�A%U�~�G
髯@�U�<�.��e�����;�[�w�\OTf!�s'�pھ�FG�Iy r%�D
�!_��T����nd�Z~z��s	����1ғ;�j�0�J��oE�;KD�������0jD�𻉆L#���} ���yP�AZ��F�"�v�����A�g����� in�(�E�?�Cx�߸���^�a�����8��LLޢ�T��ؘSg4�wM����sޝy�)�&�=I ]�{�7;v�?>�ܼ����B;��wK�2�I��Q�����B)�iX֌��-B�\q�(nC�!uY�G�E���	��(�y.�M�P�O<���́_�_�ᣯ׆R��c�[��^E�n�"]�Ql�[$����ⷄ��Z�%R�~å}��x�B��������N��C�7��)�ܳ�na����SE�5҉F��%ʱ����+)g��HX~�{����_Y	���i�!f$k�n����X`�e��Y�I�F�yu}�5@}��2�IF�+u��|7���e��Mڽۄ��7�b�����������ӿ�RN���Z��H����z$d���>��D��+�3ꬖ�N8��"��J1��O4.	�i��+\Ss���Hve3���\9Cp���*�[�����V���>�c���k/������[���LY\ {�0p�%�q4��e �z���=�{����|wn��I�	~���|���q�I������z�+?A�G��;w��3ﲥ�P���M�4�Z��"�Dd*�������nQ��J���Bn�[X=���z�Nk�����1� �l�.[N8ikM0((��f�;���:��'�0��i.˘$�/��=��覂
��΅�����������i10���o���*���4��(���R�
���]Q�Kt��}��h#9������X�"��v��ڎKR+V|��`13�#�R�j~��~�p�,��>���$<'�`u��T�5��.�	8��DRl?�u����[��)�l��x��;&�.+V�����n��ל8�o����Ӏ���CG�u4p���r�ś��]�P���K\�Iv��î��F	�9$��P�����-�KJ���N�<V���Ú�%�f7�sc,�Pm<֮�|	}��t�1e�(��;���4YI�]�~���%T�ش��y\B�U\�!t���VЍ��<��T���_l$[�IP���2�Q!��+z��8�c��Һ$�"�(ʕ��7�M�K⸆���ܷ�9+8��Me�����p��1��4�����nC�&9�Ÿ��R��Am�5����C:�院��
�eZ�jF�xj���+�숵+�3�AZ&�uh�ϑ=]5��%��R2"��uV��e�i��C!�^�\vۀT8w�Ei+Wa˟��.�8~��D^ҧ.������t�}[*�s��U�V33�$�P~�XA׺U+�lu�C��K�t�)�Zz�5m${�0�ٳ��ŵ/#�!���Ӧ�����9�:�#)�&'r�� [e$�隶��N����ay�z��C�|�\.��+�-���X���"�O#* ;I���pk��dw�LsO�d�:L�#A�����Q��g��x�k���Ƿ�Ò����X�_�6�t;6��_hr�`Uܺ�a*��;Wdx��ab�����w����0�:���Ox7�$�>� ��'���V���E�k������X���	~��2Yg�LW7K�c';��Jq�-5r쭄}�L\w�J�����r4�\67�ϼ6��E���F�(�=I+A�cn����Qv��g��Z~ZK3*(G��z��\�
0I��WG�t�0)��?\��;�������N��'ʭ�q��DC�D�!�x�WdI��\��>���N�E�x��@B��m����~���Q�ݠ��Y�����
���C5R�����X��Q�葑��K���7����!��w��B �{.�	�?����L�� t���q�i�� Ȗ;J�h� 4�Q��P�җ�F��P��4��s�l��Ei&����s��`?BoN�%�o�Q�Ή�81x��%��]72�6�PQ���_E9�0�c��:�ۚC��\��^�4�����a��d�.���1�rS_
����v�p�ˑ�
�}����ܛ��t1)N˖��S�>�x�<g����7�5o����2�����w�^D+KfY���
(g�����J����r�n��Q�EK��q.v5e	�F@^�2�F�Bꩆ�צf��w$��,�|}D�t�P��U�{��e�I��W��C��A�@]�k�#i���p����s����oz�	{��X�,xK.t�{�	V���� �� ��v�nPW�"�k���v$OԤ���J�7�}�yǍ|�PK�(ra#R�:�hh�ڝޏ�f3D�|!�9%IC��{�i��z��ti��xu�Og��kk*���Ě78��j�UEԞ���*6!�]x۹QK��z4K;�f�x����G2���eO�O��e�����$��Y��힬%h�&w `L
���S�}��u�'o�]��L臑�)Q�T����I��������8���A'.����2��Z���④�qWtZ�~ޞ�ZG[ۅ�kc�u��X�ش�#e`�@g�"Qį�?�{P�1��V��Oc���}��<�����jw7)�HEjנ�5J�,1�����2���:��$3�� �z�(bL��4��u7�ڬ	aV����@!jdHѮܖ�c�Ë�%8�)����r�D3"E�UZ�*�1h���v��� mj���m<K �''���Eq�|��Wɝo�ёz�4p:d�-���ٵ���)ЅN��.(A��/ɭR���'��B��,�7ʮ�e��O�����ɫ�p'��6�:�1渪�����q�I�����k{��Es�dK�8��$�{W�9��������8���NH�yi5�;R�|)��C&Zd��0�M�p�g��#{�#�.N�*��)��.��q$=�2$���j~s,s�ԕ�n'��~�X�wu�V9
����v Պ�c>��v��ty&�%Ȓ�$�7oQ�~�'*��V�W�XZXp��wz�A勒�*�N��ߝ8�B}�5�/� X���s�,�6IY-%i����h/$��uZ�c?�5�0i4��*%���>uu�Պ���Ԍ�R�Y4�M$s�YUkQ���)�e�h(����b�r��x/1 }��%āXFY�䧯�5��C;;mA.���u{�,�/#�֎T�<7�=��K�*ϴZ�<y�GhB8.���[��Ŵ�in�������1�Q�(K��z�"e,��2�7�
g���[z�n�1;1����P/�x4�f��<B�'zS:A,�!i�g�PM��
���6���W�뉜����E�ep��M�<h�1qR�bӟ �����$�M��M�o?E� mJ��6�{���Zs�m��y��e�>�xm���#P� ����0zlż��@fjl�ٕ�i�G�� �KZC!j�8(��Z�r���(d̈́׏���吉mb/U�K��Q�U��O~3���Uk}���z�DQ��x�#��smC��4�Gdy��n$����]b5w���^�{l:u��embޟ^KB�tƢ�%Č��Y�>1�;t,�x��۟kx�	�V�mn��d�J��WzV�@���v,"�`cQũ���RG��`���hg���&B�(�q��hJT��,5.�`m�����MP �W����;�??]<��U+�?t+�F��b/�Z� �/��ۥ��a��l�?SZ���>3Ǿ�����N�+�J�\;����5֎P��� -|�����ù�9���4�e_:w�%�x�c�^���S�����Z�F��FR�\㌎�E7�-�o,��%[<�o:�5��$n��M�ڿ�*՛e�� |�r�%Oʜ�{�aU�S'&���52��Xƭy;�R�!	?ӓ_)]�9��x�nd	#}P��.#�x�z�H��ʒ/
:�3��|��%)��(ӧ��m�{��y��N��M��H�wh�|�K�୯2��5�>���F� �p������L�56�8[���Y����I}b�A���,��)�T���`�z.3X"`�i_`V�+	��2�i�Z)Ό�Ӑ���A���Leu��`��D1_Z,EhУ��`�u�ɣ &�J&�!�̇�{ߥ�y�hL6T%4H�[�9`�8��^4��#Ow3^�~��@G= � ��g�-�*m�ش���F�B�Ǝ�p5&�S��?c�,0@�TU,�$]�b�J�CH;�2}�n<E�*<VW��f��"7���
h�VϽ�ƞ8�xz;~�&�rC�����%���+8}c����C+2Ⱈ���Oh���0ڑ�>Fu!��<�Ue�*��ؿ.���xTda�'Ē�YC�G��ݝ�oF��6âS<װ�Ti�8�K���w�X���eTG�ap@�����jt o����Ol~��l�@��n��Ń��[ؠ2 l<"���f�^���m�SXw*_1�&��N|'�WG�e�w``a�r��G�2|���ֳ�f�q���Lգ�jyR��Z��c^�&�Ѷ2b.�hg`�R3E�R�����h�Co]t�����(VS~g��pO�y�̴= Gw���e��gddp4N' �l[l�u�Y��#ډ�/���Q�طN#y^pB�VB����r+�Z�脿��>d��9JN���`�@zW���ӭ_�-��`4>��x/*�pP���gΟ��?Ёt�RF�@9P�{�����%��+�r���qW�p�7@K��fpK��p����gL��Fu/�*Do��P�j	>��� /���� mD��l��9{�'���%:f]i�Rݠ���r�I�3
N�"�f. �!XxFn���6V)¢H�`PN��7.��G���x�ž����/1���4����,�#��S��F`Z�ZW�m	/�V�ã�Vq4��/pA�$����P|�b���� ��I�9���$�T�C}+z*��w���,}�P��t�Sȸ�sz���bǝQn�
� >��N96"M�U���iA)x6
^0 �� �:u#��K��9 u�f�I��(�m+�(��T|��b'����0��g\��(kϩ@B�����R����@��`�������S� :{X�WW�s�Ke���2нT7���8�ͨ-ǈ@KHQ�� ��W:� B�?�M,����A�b�=f�d�kx�z��7U���1��#)�^2%���j;�}<��QP#P�d�͊=���w�e��`ڝ�M�ŕC5�FÇp�B �x�T�B<�䗙;y�,s1@��|L��5X"�6_u�7�{O�qV�n�0'�P���kdK��0J8�^�M'*���Y5�?�Pk|�&@��jzA_w�c�M�K��);J��ް��"��EMh�����Uany�Jn�>w#7�tjV�[k�"�2Πn�F��}sU]�-����~�1[.nҜXl�;޽�B��aN%kJy��6�A�].o`D�%AZ���4T�}��+1���t���b6��]O��t���<}��/Y��.sxa�v��9��g�s��^o��G#��O�%lm��m��f�5LպD<*�-
�YW`Q��S���#Iŏ(~Ԧ��*�u8�F�; �'���a���#�^,��)����Ƙ�� �)���$�SpO]�c���Iש��%Cy[�>�EнC.[?}���L���}�$\��>1P����M3�rB�#L�\�{�g�1�)9���X�3
̜d��pժʸ���w��6�cH�ȅȍr<����0ywc]Q�-`�Z+�~�(.Xa�-�'6�ac�1a~��o.O#ָy�l{^�g�^3Y�ǚ-Bә� ��K���rO�J~��.���4�W��2�hB>I���瑶���U���b����@]Y�A�h~��_���Ҝ+
V�cT����Zl��~�����l�J�3���B�}uv���쇇�B���Έ.Im���?D���"���x���y��C�� <�O]W(r*��v�R�ނ�eG��6L#d�/�����g:T�ͬ�ð��i�<(���DQ`*�	p��:�Q�N�|��"l���|�WE��^���$�\)*��s������&
'��@���CƜ�Բ�/癛���>�ڂ�qu�Ϫ��z6m#���i� ҕ�ۖ��,r�t� �ih�,�D�'ȐX�iQ�q,Sח).C.���:�<f�y�W��F^��G�BD<��������/�>:�Q��� �p���zd%�K���a(b�+?MF#�"���\-C�������EQ���7���q��d�`!F��Q��|w�e6��VY�ژ�eվ͹�v�������O�<!S�
���c�v;TZx/��uVy�0�(�Ha+=_\Ӎ�޿���jc��W��W�;>9���a�� ��9cEC��zWs���İ:ދ���)�꽃��5� �n^������;�fy�b�CU
�NbBP�����,y��ykF)��9����G��#��qtA��AJ-R��a�j��1�U�G������ŎvI+[�X�pok�#��f�[:����",(Tv"�<%D��ME����y�Y��1[��5�bP�	���}١��(�H���F��S�����"�n
؍�E��	0�`T��_���ל�g��ғi�׾vej�\��+�z����m�jmǖ nZ�骒|�ÎR_i�k;E��EV�e`o�p�+�%M�U��h^�ʞ�b���H�Y9W�����af2M�Y<�'�(����D����{����J˻p��##�o�H,,��R�W�C�t�	�O����Gē��3WUKjTe���ћ���ǓF���n��b��#v9��p�����huF-h����f�[i?�3Ta+�LޭS�݉�=��i����Od~Y!��*�j�����w<���$b�£'�M|R��%g�A�/�>�'AF֝�%���A|F���Y���a6���q���١a=�	"��*#
4�LA\$b����?C�'|D"p���oci,��
35� A>w�u��1��0ּ�¾�ʓ���ف���I\�.��Ե���tM�,))�����ʔ:a6ui���Nkᶓ�p�*�|��qF�L;M�S�$Z��q��xc��,��^��e�����\���sB�����p\;���t�fD&zU�#�[���K%�i6�(�)�	���r:X�a���Z�-
SL� �j �N�k\��n�����-��qޱJ���:��}�m 

2� c�ye��DI�(��o�Y�*���龿�W0Ӿ9v�	B�{�A�i9�6U��t�,��|�Z�Pk�:��m���z��\��M�M�7ɬ�+^��%�+���C�L��*<7��_�ڏ�H���������8�w��Z�z��Y��W�^��@�9?!s���_��@Q���c�����]���	-�t�G���k���U��U"�,IWQl!E�o"dT��6 |#s��Vڙ�Zo���;N�s?�:Y��� 1������{��;�sR��k�y���ʩ%���N̬��^kң�(�|�����G���ppB؟I�A�S�@��L>�-�Tż����^��)s�B9���3V`�㸻1	#l�10m�b�8�/$��?���=������\�#&t[�|^ٚ�)�
U�񥐃]�;�sUlN����p�pvq�/y	#�bl�`�<ۼ�.���gj���='=ɞ�R;�ؘER�)��.@�޳Y�Z�M�%�ϓ���4%t������MIM!�!����;�R����8��/K.��-ߜr�w�e!n���vP)�gi���</'�C4�bDl����'�}I��+5������R��1+�9����QN�tTX���h�"�=�v �Ԓ2<�{N�c���dH�6��RzD���7zZ$��p���F��7���q�d%PI�Z��M�����D�k�k/�!٘�C�Z��{���5���Є���n�B�����(���g�.O����ӆ�?ԳGv�-�3H�%z��=z�.m^Jܰb����m��\�c�eZ�&��h�:#�G;�i	�y���CH4CժM�j]�Ƶ���zK<��� 1�z���`��X�B�>���%�/����M�q�o��L��|��S$uG��j�����g�@&��$^c�%�2�q�t�cr��b��9��M��]�_�Lw��� �/��ǂ�?N���I{��)נiҵ����&���+F<����h �M��A����A$@0s�񇣆4�u���:�B�5��C�^�� �K�	m��)Z�}�<�h�/@)8Z�@ٹ��aпk�A$�a�|�pP�R^��\d�o����@\����^��ک,`�L��M�,C]���ZԷCX�s�Ų�͜#i<��.��k�Aݍ�łh�u$ڀ{3񬓸����ά=��T����7J�2c;LH�RHq��	�"��;���53�%�l���P/��7���9�)mg� �J=����@��k���k���_ck��
��A}&���c��ı��hJ[�EkZ����i_�0 �L>U���Z�Ӷ�z��)��Au_#�.�B�b{u~�v1�&����ї���@)/w�$�>JD�ߓ�$p4�/C�Z�o��=�jt���o�ξė��.���*�0����@r#�m�n>$�Q��AR�i��Z:BfN�Z4�~�\���2��c!ZԵvp�r݈� ���D���oH^�%��ţn�T�z1�"^d�:-<%�=�54����P�����%��b�&:]�ޛS���b62r��8��%dh�6�  H��Q(r� !�v�-g�������cT�m�����}6ז��U�/�����Y�����1�<��Q{8��y9�8��{��S��1z�%���#v����ZN_�}�
q�A�����d��W�g^���mz�7� �׉w>!�����XB����dM�W���� !֣`��4h�g;��0��a��?m���s'��Z��,K�G��O���aKj���0�Q��J��񕣁�rQc8hmͣ�6lQR�����1���+n~�c����AKkk�M�SL9A�2]����8�C}��2E�]���	��7���}��-��YQ���]Ma<����S~��� >a��w6*nx�FkI�Xl����OB��g�)��BWs=Z�"���H�H�<q��c۳����@&�RZɢ���%gg�oTĳPX���}���K��}R�
����� �� �]��3�+r�����)!�`�AY��]�0��;�|��aל�ӷ���f���+����l�9s4Pvm�ףZ�ѳg�VW����<G�*Ҙ|8�ѝ7�#R��c������P��!IT�S��G�\D�:ѭcr��p�S��U�z�c����gaE@}!��YSXg�D	��>gd z�U����z�02��g(�Kbq�����V#{��Cw�n�ݖ��5���.n
�ߗQiuJ�n�zq�-���l�m2�⨨����L_�,cpWݟ/�I{�����Z�F�>|jyq��~�	��:Nu��h�Hߡ���k �2��h��V y�B�JO���=�I�h�̿�d��P[�6����R�c���`��_��4^C�~S	I�eW��~�ɣ("�f4��4!����_~fI��4�+�Ҷm��=r��S�Ӳ�.�����ϾK7s����-1$jS2�:UjĐ�W'�4��`	r~��ݪ͙PS!��Iܣ�.�����YI�L�z�\�
�!M.�д�mF�6U
����I���ɬ���<׆T�j�8�8�'�<Ex�1������+
��:;�{��L���4{qu��^7.�׫�$�uN"�qS�%1�I�C��t=�h@6��0T_B�+ׅ��[���5&(�'�l0G�d�p���3�[P
�A'�S�{R��*��߇Ds����)�@��Q� 1�B��@��n��<�4�����M�'l|/O�I�����W��Cz	�_ÇY��=��^D�X����5��|��f[�^�DM�b��9��t<�V�����VR���<(���$�Us���~�`;�f�L�nv=��[�'��������_ߺD���
�6�tR���y�^IV=�R��O:�<�F+Q��eeiD�����0	�F����|�1oZyT�p�e?�iW~�z8�<���˯�#��	��>~��\=���(������p\<ͻ���7d7m��,�����b�f�ta�Ī_��@G6X�r���'��r$;l�������D�0%��s�h	u���淭/�$��m�\���Z���e��d��{�'(�����Д���G�TU{���G�GT����Q-Ǣ�����#(������M��|�׆�%oǃ!�h�[�>�,q��Ї+�e��(�q�7H#��	�@�<��'->��w��v���w�@KU��D�0����lХ�0A �rK�Ѥp�꣋<C���N(�4N⦕��Wv5�>N����"��*ȡ�Ι}D;���9B�^�����r4�y�yjއ*n��Qݵ�-0ȖԆ>K/=��w�c�E�Mx����ߣ?M��5OQq1�O4�	|�"c_�'��<1�x�]��-�4���%�c���B�ۄ�W�|,!���Ooԥ�|6٫��-Z��,�Lf��ǤjR���4�05��:g�b)k�y[->̀"��m�E�����CNd%��<H���e�;O�Ѝ޳�!���(��6���MB^om |^[SΩ��~���X3���������&��|CP��P�.p��!j2�a{���S����	���;$�H��=�<��sw��K0�]�dg��fV�/� -��[pQPa�@����nZ;ɺ>�6ݪ{��B��V
@�X��Aq]]0��@��E֢ &-F�(�ź�"�:[����u�)¯=�lV���x�X:O]V!�Նޙ����[FN4qs�9%q>j�f�fv&�VōPs�?�>�k��3�cI�s�$M���,����|<�xʬ��ΣXQ��&y�kl.�HW��o���<��2��+2Y�j����Y�j��E�����_�-~ق�1�j�aJ����� X�e�_n(��$�t�������-��m�ʃX�*�R��T�A�J�-�m�W��@F����{�#P�J�?� �nQ��a��v���<�oH��lu��T�5+^�DC���^���Ԙ��������e/��PRcJ�tx��u6�u�*���KR
�y8�v�.��5�F.��T,h� �&��U�{�L#1�R~�.S�����R#�vc��֘P@!�}����袥�UU�e�L2~F�G��^	�\a��e��A�ڻ������D>� ��H���c��$�I�}:~���s�i��]lX������;�O��]���6?Pk�z�e�͆��Ǻϵ���$ Q�<ʙwQ$h���E�i�֨�׵dsd�Εۥ�\F�����4C[��)��A���1������ѿ�bWJE0Yw�^-h��R�&�Ag�������3l�10����p���T�ŝ?9m��os�t��ƞl-E_Y�������C�!m�����ЯKy���qcq3X�g